magic
tech scmos
timestamp 1700564293
<< nwell >>
rect 462 557 498 589
rect 518 557 554 589
rect 573 548 609 580
rect 637 557 673 589
rect 693 557 729 589
rect 748 548 784 580
rect 812 557 848 589
rect 868 557 904 589
rect 923 548 959 580
rect 987 557 1023 589
rect 1043 557 1079 589
rect 1098 548 1134 580
rect 1165 557 1201 589
rect 1221 557 1257 589
rect 1276 548 1312 580
rect 1335 557 1371 589
rect 1391 557 1427 589
rect 1446 548 1482 580
rect 1505 557 1541 589
rect 1561 557 1597 589
rect 1616 548 1652 580
rect 1675 557 1711 589
rect 1731 557 1767 589
rect 1786 548 1822 580
rect 462 406 498 438
rect 518 406 554 438
rect 573 397 609 429
rect 637 406 673 438
rect 693 406 729 438
rect 748 397 784 429
rect 812 406 848 438
rect 868 406 904 438
rect 923 397 959 429
rect 987 406 1023 438
rect 1043 406 1079 438
rect 1098 397 1134 429
rect 2469 348 2505 380
rect 2532 348 2568 380
rect 2647 348 2683 380
rect 2710 348 2746 380
rect 2802 348 2838 380
rect 2865 348 2901 380
rect 2958 348 2994 380
rect 3021 348 3057 380
rect 2353 312 2389 344
rect 616 233 652 265
rect 672 233 708 265
rect 727 224 763 256
rect 786 233 822 265
rect 842 233 878 265
rect 897 224 933 256
rect 1160 246 1196 278
rect 1216 246 1252 278
rect 1271 237 1307 269
rect 1335 246 1371 278
rect 1391 246 1427 278
rect 1446 237 1482 269
rect 1510 246 1546 278
rect 1566 246 1602 278
rect 1621 237 1657 269
rect 1685 246 1721 278
rect 1741 246 1777 278
rect 1796 237 1832 269
rect 2533 263 2569 295
rect 2711 263 2747 295
rect 2866 263 2902 295
rect 3022 263 3058 295
rect 558 177 594 209
rect 2265 135 2301 167
rect 2321 135 2357 167
rect 616 95 652 127
rect 672 95 708 127
rect 727 86 763 118
rect 786 95 822 127
rect 842 95 878 127
rect 897 86 933 118
rect 1007 99 1043 131
rect 1160 95 1196 127
rect 1216 95 1252 127
rect 1271 86 1307 118
rect 1335 95 1371 127
rect 1391 95 1427 127
rect 1446 86 1482 118
rect 1510 95 1546 127
rect 1566 95 1602 127
rect 1621 86 1657 118
rect 1685 95 1721 127
rect 1741 95 1777 127
rect 2376 126 2412 158
rect 2447 135 2483 167
rect 2503 135 2539 167
rect 2558 126 2594 158
rect 2640 139 2676 171
rect 2787 135 2823 167
rect 2843 135 2879 167
rect 2898 126 2934 158
rect 2969 135 3005 167
rect 3025 135 3061 167
rect 3080 126 3116 158
rect 3162 139 3198 171
rect 1796 86 1832 118
rect 2640 93 2676 125
rect 2728 86 2764 118
rect 3162 93 3198 125
rect 3250 86 3286 118
rect 558 39 594 71
rect 1007 53 1043 85
rect 1095 46 1131 78
rect 2324 -3 2360 29
rect 2387 -3 2423 29
rect 2635 0 2671 32
rect 2698 0 2734 32
rect 2846 -3 2882 29
rect 2909 -3 2945 29
rect 3157 0 3193 32
rect 3220 0 3256 32
rect 2324 -85 2360 -53
rect 2388 -88 2424 -56
rect 2635 -82 2671 -50
rect 2699 -85 2735 -53
rect 2846 -85 2882 -53
rect 2910 -88 2946 -56
rect 3157 -82 3193 -50
rect 3221 -85 3257 -53
rect 505 -151 541 -119
rect 561 -151 597 -119
rect 616 -160 652 -128
rect 680 -151 716 -119
rect 736 -151 772 -119
rect 791 -160 827 -128
rect 855 -151 891 -119
rect 911 -151 947 -119
rect 966 -160 1002 -128
rect 1030 -151 1066 -119
rect 1086 -151 1122 -119
rect 1141 -160 1177 -128
rect 2265 -251 2301 -219
rect 2321 -251 2357 -219
rect 2376 -260 2412 -228
rect 2447 -251 2483 -219
rect 2503 -251 2539 -219
rect 2558 -260 2594 -228
rect 2640 -247 2676 -215
rect 2787 -251 2823 -219
rect 2843 -251 2879 -219
rect 2898 -260 2934 -228
rect 2969 -251 3005 -219
rect 3025 -251 3061 -219
rect 3080 -260 3116 -228
rect 3162 -247 3198 -215
rect 505 -302 541 -270
rect 561 -302 597 -270
rect 616 -311 652 -279
rect 680 -302 716 -270
rect 736 -302 772 -270
rect 791 -311 827 -279
rect 855 -302 891 -270
rect 911 -302 947 -270
rect 966 -311 1002 -279
rect 1030 -302 1066 -270
rect 1086 -302 1122 -270
rect 1141 -311 1177 -279
rect 2640 -293 2676 -261
rect 2728 -300 2764 -268
rect 3162 -293 3198 -261
rect 3250 -300 3286 -268
rect 2324 -389 2360 -357
rect 2387 -389 2423 -357
rect 2635 -386 2671 -354
rect 2698 -386 2734 -354
rect 2846 -389 2882 -357
rect 2909 -389 2945 -357
rect 3157 -386 3193 -354
rect 3220 -386 3256 -354
rect 628 -477 664 -445
rect 691 -477 727 -445
rect 769 -477 805 -445
rect 832 -477 868 -445
rect 913 -477 949 -445
rect 969 -477 1005 -445
rect 1025 -477 1061 -445
rect 1081 -477 1117 -445
rect 1133 -486 1169 -454
rect 2324 -471 2360 -439
rect 2388 -474 2424 -442
rect 2635 -468 2671 -436
rect 2699 -471 2735 -439
rect 2846 -471 2882 -439
rect 2910 -474 2946 -442
rect 3157 -468 3193 -436
rect 3221 -471 3257 -439
rect 628 -559 664 -527
rect 692 -562 728 -530
rect 769 -559 805 -527
rect 833 -562 869 -530
rect 1230 -542 1266 -510
rect 1286 -542 1322 -510
rect 1342 -542 1378 -510
rect 1398 -542 1434 -510
rect 1453 -542 1489 -510
rect 1592 -613 1628 -581
rect 1648 -613 1684 -581
rect 1703 -622 1739 -590
rect 1762 -613 1798 -581
rect 1818 -613 1854 -581
rect 1873 -622 1909 -590
rect 1932 -613 1968 -581
rect 1988 -613 2024 -581
rect 2043 -622 2079 -590
rect 2102 -613 2138 -581
rect 2158 -613 2194 -581
rect 2213 -622 2249 -590
rect 628 -658 664 -626
rect 691 -658 727 -626
rect 769 -658 805 -626
rect 832 -658 868 -626
rect 943 -694 979 -662
rect 999 -694 1035 -662
rect 1097 -694 1133 -662
rect 628 -740 664 -708
rect 692 -743 728 -711
rect 769 -740 805 -708
rect 833 -743 869 -711
rect 1097 -740 1133 -708
rect 628 -839 664 -807
rect 684 -839 720 -807
rect 740 -839 776 -807
rect 836 -838 872 -806
rect 892 -838 928 -806
rect 948 -838 984 -806
rect 1004 -838 1040 -806
rect 1128 -838 1164 -806
rect 1184 -838 1220 -806
rect 1240 -838 1276 -806
rect 1296 -838 1332 -806
rect 1410 -916 1446 -884
rect 1466 -916 1502 -884
rect 1521 -925 1557 -893
<< ntransistor >>
rect 505 511 509 531
rect 589 518 593 538
rect 680 511 684 531
rect 764 518 768 538
rect 855 511 859 531
rect 939 518 943 538
rect 1030 511 1034 531
rect 1114 518 1118 538
rect 1208 511 1212 531
rect 1292 518 1296 538
rect 1378 511 1382 531
rect 1462 518 1466 538
rect 1548 511 1552 531
rect 1632 518 1636 538
rect 1718 511 1722 531
rect 1802 518 1806 538
rect 505 471 509 491
rect 680 471 684 491
rect 855 471 859 491
rect 1030 471 1034 491
rect 1208 471 1212 491
rect 1378 471 1382 491
rect 1548 471 1552 491
rect 1718 471 1722 491
rect 505 360 509 380
rect 589 367 593 387
rect 680 360 684 380
rect 764 367 768 387
rect 855 360 859 380
rect 939 367 943 387
rect 1030 360 1034 380
rect 1114 367 1118 387
rect 505 320 509 340
rect 680 320 684 340
rect 855 320 859 340
rect 1030 320 1034 340
rect 2485 318 2489 338
rect 2564 309 2568 329
rect 2663 318 2667 338
rect 2742 309 2746 329
rect 2818 318 2822 338
rect 2897 309 2901 329
rect 2974 318 2978 338
rect 3053 309 3057 329
rect 2369 282 2373 302
rect 659 187 663 207
rect 743 194 747 214
rect 829 187 833 207
rect 913 194 917 214
rect 1203 200 1207 220
rect 1287 207 1291 227
rect 1378 200 1382 220
rect 1462 207 1466 227
rect 1553 200 1557 220
rect 1637 207 1641 227
rect 1728 200 1732 220
rect 1812 207 1816 227
rect 2565 224 2569 244
rect 2743 224 2747 244
rect 2898 224 2902 244
rect 3054 224 3058 244
rect 574 147 578 167
rect 659 147 663 167
rect 829 147 833 167
rect 1203 160 1207 180
rect 1378 160 1382 180
rect 1553 160 1557 180
rect 1728 160 1732 180
rect 2308 89 2312 109
rect 2392 96 2396 116
rect 2490 89 2494 109
rect 2574 96 2578 116
rect 2830 89 2834 109
rect 2914 96 2918 116
rect 3012 89 3016 109
rect 3096 96 3100 116
rect 659 49 663 69
rect 743 56 747 76
rect 829 49 833 69
rect 913 56 917 76
rect 1203 49 1207 69
rect 1287 56 1291 76
rect 1378 49 1382 69
rect 1462 56 1466 76
rect 1553 49 1557 69
rect 1637 56 1641 76
rect 1728 49 1732 69
rect 1812 56 1816 76
rect 2308 49 2312 69
rect 2490 49 2494 69
rect 2646 53 2650 73
rect 2697 53 2701 73
rect 2744 56 2748 76
rect 2830 49 2834 69
rect 3012 49 3016 69
rect 3168 53 3172 73
rect 3219 53 3223 73
rect 3266 56 3270 76
rect 574 9 578 29
rect 659 9 663 29
rect 829 9 833 29
rect 1013 13 1017 33
rect 1064 13 1068 33
rect 1111 16 1115 36
rect 1203 9 1207 29
rect 1378 9 1382 29
rect 1553 9 1557 29
rect 1728 9 1732 29
rect 2340 -33 2344 -13
rect 2419 -42 2423 -22
rect 2651 -30 2655 -10
rect 2730 -39 2734 -19
rect 2862 -33 2866 -13
rect 2941 -42 2945 -22
rect 3173 -30 3177 -10
rect 3252 -39 3256 -19
rect 2340 -115 2344 -95
rect 2420 -127 2424 -107
rect 2651 -112 2655 -92
rect 2731 -124 2735 -104
rect 2862 -115 2866 -95
rect 2942 -127 2946 -107
rect 3173 -112 3177 -92
rect 3253 -124 3257 -104
rect 548 -197 552 -177
rect 632 -190 636 -170
rect 723 -197 727 -177
rect 807 -190 811 -170
rect 898 -197 902 -177
rect 982 -190 986 -170
rect 1073 -197 1077 -177
rect 1157 -190 1161 -170
rect 548 -237 552 -217
rect 723 -237 727 -217
rect 898 -237 902 -217
rect 1073 -237 1077 -217
rect 2308 -297 2312 -277
rect 2392 -290 2396 -270
rect 2490 -297 2494 -277
rect 2574 -290 2578 -270
rect 2830 -297 2834 -277
rect 2914 -290 2918 -270
rect 3012 -297 3016 -277
rect 3096 -290 3100 -270
rect 548 -348 552 -328
rect 632 -341 636 -321
rect 723 -348 727 -328
rect 807 -341 811 -321
rect 898 -348 902 -328
rect 982 -341 986 -321
rect 1073 -348 1077 -328
rect 1157 -341 1161 -321
rect 2308 -337 2312 -317
rect 2490 -337 2494 -317
rect 2646 -333 2650 -313
rect 2697 -333 2701 -313
rect 2744 -330 2748 -310
rect 2830 -337 2834 -317
rect 3012 -337 3016 -317
rect 3168 -333 3172 -313
rect 3219 -333 3223 -313
rect 3266 -330 3270 -310
rect 548 -388 552 -368
rect 723 -388 727 -368
rect 898 -388 902 -368
rect 1073 -388 1077 -368
rect 2340 -419 2344 -399
rect 2419 -428 2423 -408
rect 2651 -416 2655 -396
rect 2730 -425 2734 -405
rect 2862 -419 2866 -399
rect 2941 -428 2945 -408
rect 3173 -416 3177 -396
rect 3252 -425 3256 -405
rect 644 -507 648 -487
rect 723 -516 727 -496
rect 785 -507 789 -487
rect 864 -516 868 -496
rect 956 -523 960 -503
rect 1149 -516 1153 -496
rect 2340 -501 2344 -481
rect 2420 -513 2424 -493
rect 2651 -498 2655 -478
rect 2731 -510 2735 -490
rect 2862 -501 2866 -481
rect 2942 -513 2946 -493
rect 3173 -498 3177 -478
rect 3253 -510 3257 -490
rect 956 -563 960 -543
rect 644 -589 648 -569
rect 724 -601 728 -581
rect 785 -589 789 -569
rect 865 -601 869 -581
rect 956 -603 960 -583
rect 1273 -588 1277 -568
rect 956 -642 960 -622
rect 1273 -628 1277 -608
rect 1273 -668 1277 -648
rect 1635 -659 1639 -639
rect 1719 -652 1723 -632
rect 1805 -659 1809 -639
rect 1889 -652 1893 -632
rect 1975 -659 1979 -639
rect 2059 -652 2063 -632
rect 2145 -659 2149 -639
rect 2229 -652 2233 -632
rect 644 -688 648 -668
rect 723 -697 727 -677
rect 785 -688 789 -668
rect 864 -697 868 -677
rect 1273 -707 1277 -687
rect 1635 -699 1639 -679
rect 1805 -699 1809 -679
rect 1975 -699 1979 -679
rect 2145 -699 2149 -679
rect 986 -740 990 -720
rect 1273 -746 1277 -726
rect 644 -770 648 -750
rect 724 -782 728 -762
rect 785 -770 789 -750
rect 865 -782 869 -762
rect 986 -780 990 -760
rect 1103 -780 1107 -760
rect 1154 -780 1158 -760
rect 671 -885 675 -865
rect 879 -884 883 -864
rect 1171 -884 1175 -864
rect 671 -925 675 -905
rect 879 -924 883 -904
rect 1171 -924 1175 -904
rect 671 -965 675 -945
rect 879 -964 883 -944
rect 1171 -964 1175 -944
rect 1453 -962 1457 -942
rect 1537 -955 1541 -935
rect 879 -1003 883 -983
rect 1171 -1003 1175 -983
rect 1453 -1002 1457 -982
<< ptransistor >>
rect 479 563 481 583
rect 535 563 537 583
rect 590 554 592 574
rect 654 563 656 583
rect 710 563 712 583
rect 765 554 767 574
rect 829 563 831 583
rect 885 563 887 583
rect 940 554 942 574
rect 1004 563 1006 583
rect 1060 563 1062 583
rect 1115 554 1117 574
rect 1182 563 1184 583
rect 1238 563 1240 583
rect 1293 554 1295 574
rect 1352 563 1354 583
rect 1408 563 1410 583
rect 1463 554 1465 574
rect 1522 563 1524 583
rect 1578 563 1580 583
rect 1633 554 1635 574
rect 1692 563 1694 583
rect 1748 563 1750 583
rect 1803 554 1805 574
rect 479 412 481 432
rect 535 412 537 432
rect 590 403 592 423
rect 654 412 656 432
rect 710 412 712 432
rect 765 403 767 423
rect 829 412 831 432
rect 885 412 887 432
rect 940 403 942 423
rect 1004 412 1006 432
rect 1060 412 1062 432
rect 1115 403 1117 423
rect 2486 354 2488 374
rect 2549 354 2551 374
rect 2664 354 2666 374
rect 2727 354 2729 374
rect 2819 354 2821 374
rect 2882 354 2884 374
rect 2975 354 2977 374
rect 3038 354 3040 374
rect 2370 318 2372 338
rect 633 239 635 259
rect 689 239 691 259
rect 744 230 746 250
rect 803 239 805 259
rect 859 239 861 259
rect 1177 252 1179 272
rect 1233 252 1235 272
rect 914 230 916 250
rect 1288 243 1290 263
rect 1352 252 1354 272
rect 1408 252 1410 272
rect 1463 243 1465 263
rect 1527 252 1529 272
rect 1583 252 1585 272
rect 1638 243 1640 263
rect 1702 252 1704 272
rect 1758 252 1760 272
rect 2550 269 2552 289
rect 2728 269 2730 289
rect 2883 269 2885 289
rect 3039 269 3041 289
rect 1813 243 1815 263
rect 575 183 577 203
rect 2282 141 2284 161
rect 2338 141 2340 161
rect 2393 132 2395 152
rect 2464 141 2466 161
rect 2520 141 2522 161
rect 2575 132 2577 152
rect 2657 145 2659 165
rect 2804 141 2806 161
rect 2860 141 2862 161
rect 2915 132 2917 152
rect 2986 141 2988 161
rect 3042 141 3044 161
rect 3097 132 3099 152
rect 3179 145 3181 165
rect 633 101 635 121
rect 689 101 691 121
rect 744 92 746 112
rect 803 101 805 121
rect 859 101 861 121
rect 914 92 916 112
rect 1024 105 1026 125
rect 1177 101 1179 121
rect 1233 101 1235 121
rect 1288 92 1290 112
rect 1352 101 1354 121
rect 1408 101 1410 121
rect 1463 92 1465 112
rect 1527 101 1529 121
rect 1583 101 1585 121
rect 1638 92 1640 112
rect 1702 101 1704 121
rect 1758 101 1760 121
rect 1813 92 1815 112
rect 2657 99 2659 119
rect 2745 92 2747 112
rect 3179 99 3181 119
rect 3267 92 3269 112
rect 575 45 577 65
rect 1024 59 1026 79
rect 1112 52 1114 72
rect 2341 3 2343 23
rect 2404 3 2406 23
rect 2652 6 2654 26
rect 2715 6 2717 26
rect 2863 3 2865 23
rect 2926 3 2928 23
rect 3174 6 3176 26
rect 3237 6 3239 26
rect 2341 -79 2343 -59
rect 2405 -82 2407 -62
rect 2652 -76 2654 -56
rect 2716 -79 2718 -59
rect 2863 -79 2865 -59
rect 2927 -82 2929 -62
rect 3174 -76 3176 -56
rect 3238 -79 3240 -59
rect 522 -145 524 -125
rect 578 -145 580 -125
rect 633 -154 635 -134
rect 697 -145 699 -125
rect 753 -145 755 -125
rect 808 -154 810 -134
rect 872 -145 874 -125
rect 928 -145 930 -125
rect 983 -154 985 -134
rect 1047 -145 1049 -125
rect 1103 -145 1105 -125
rect 1158 -154 1160 -134
rect 2282 -245 2284 -225
rect 2338 -245 2340 -225
rect 2393 -254 2395 -234
rect 2464 -245 2466 -225
rect 2520 -245 2522 -225
rect 2575 -254 2577 -234
rect 2657 -241 2659 -221
rect 2804 -245 2806 -225
rect 2860 -245 2862 -225
rect 2915 -254 2917 -234
rect 2986 -245 2988 -225
rect 3042 -245 3044 -225
rect 3097 -254 3099 -234
rect 3179 -241 3181 -221
rect 522 -296 524 -276
rect 578 -296 580 -276
rect 633 -305 635 -285
rect 697 -296 699 -276
rect 753 -296 755 -276
rect 808 -305 810 -285
rect 872 -296 874 -276
rect 928 -296 930 -276
rect 983 -305 985 -285
rect 1047 -296 1049 -276
rect 1103 -296 1105 -276
rect 1158 -305 1160 -285
rect 2657 -287 2659 -267
rect 2745 -294 2747 -274
rect 3179 -287 3181 -267
rect 3267 -294 3269 -274
rect 2341 -383 2343 -363
rect 2404 -383 2406 -363
rect 2652 -380 2654 -360
rect 2715 -380 2717 -360
rect 2863 -383 2865 -363
rect 2926 -383 2928 -363
rect 3174 -380 3176 -360
rect 3237 -380 3239 -360
rect 645 -471 647 -451
rect 708 -471 710 -451
rect 786 -471 788 -451
rect 849 -471 851 -451
rect 930 -471 932 -451
rect 986 -471 988 -451
rect 1042 -471 1044 -451
rect 1098 -471 1100 -451
rect 1150 -480 1152 -460
rect 2341 -465 2343 -445
rect 2405 -468 2407 -448
rect 2652 -462 2654 -442
rect 2716 -465 2718 -445
rect 2863 -465 2865 -445
rect 2927 -468 2929 -448
rect 3174 -462 3176 -442
rect 3238 -465 3240 -445
rect 645 -553 647 -533
rect 709 -556 711 -536
rect 786 -553 788 -533
rect 1247 -536 1249 -516
rect 1303 -536 1305 -516
rect 1359 -536 1361 -516
rect 1415 -536 1417 -516
rect 1470 -536 1472 -516
rect 850 -556 852 -536
rect 1609 -607 1611 -587
rect 1665 -607 1667 -587
rect 645 -652 647 -632
rect 708 -652 710 -632
rect 786 -652 788 -632
rect 849 -652 851 -632
rect 1720 -616 1722 -596
rect 1779 -607 1781 -587
rect 1835 -607 1837 -587
rect 1890 -616 1892 -596
rect 1949 -607 1951 -587
rect 2005 -607 2007 -587
rect 2060 -616 2062 -596
rect 2119 -607 2121 -587
rect 2175 -607 2177 -587
rect 2230 -616 2232 -596
rect 960 -688 962 -668
rect 1016 -688 1018 -668
rect 1114 -688 1116 -668
rect 645 -734 647 -714
rect 709 -737 711 -717
rect 786 -734 788 -714
rect 850 -737 852 -717
rect 1114 -734 1116 -714
rect 645 -833 647 -813
rect 701 -833 703 -813
rect 757 -833 759 -813
rect 853 -832 855 -812
rect 909 -832 911 -812
rect 965 -832 967 -812
rect 1021 -832 1023 -812
rect 1145 -832 1147 -812
rect 1201 -832 1203 -812
rect 1257 -832 1259 -812
rect 1313 -832 1315 -812
rect 1427 -910 1429 -890
rect 1483 -910 1485 -890
rect 1538 -919 1540 -899
<< ndiffusion >>
rect 504 511 505 531
rect 509 511 510 531
rect 588 518 589 538
rect 593 518 594 538
rect 679 511 680 531
rect 684 511 685 531
rect 763 518 764 538
rect 768 518 769 538
rect 854 511 855 531
rect 859 511 860 531
rect 938 518 939 538
rect 943 518 944 538
rect 1029 511 1030 531
rect 1034 511 1035 531
rect 1113 518 1114 538
rect 1118 518 1119 538
rect 1207 511 1208 531
rect 1212 511 1213 531
rect 1291 518 1292 538
rect 1296 518 1297 538
rect 1377 511 1378 531
rect 1382 511 1383 531
rect 1461 518 1462 538
rect 1466 518 1467 538
rect 1547 511 1548 531
rect 1552 511 1553 531
rect 1631 518 1632 538
rect 1636 518 1637 538
rect 1717 511 1718 531
rect 1722 511 1723 531
rect 1801 518 1802 538
rect 1806 518 1807 538
rect 504 471 505 491
rect 509 471 510 491
rect 679 471 680 491
rect 684 471 685 491
rect 854 471 855 491
rect 859 471 860 491
rect 1029 471 1030 491
rect 1034 471 1035 491
rect 1207 471 1208 491
rect 1212 471 1213 491
rect 1377 471 1378 491
rect 1382 471 1383 491
rect 1547 471 1548 491
rect 1552 471 1553 491
rect 1717 471 1718 491
rect 1722 471 1723 491
rect 504 360 505 380
rect 509 360 510 380
rect 588 367 589 387
rect 593 367 594 387
rect 679 360 680 380
rect 684 360 685 380
rect 763 367 764 387
rect 768 367 769 387
rect 854 360 855 380
rect 859 360 860 380
rect 938 367 939 387
rect 943 367 944 387
rect 1029 360 1030 380
rect 1034 360 1035 380
rect 1113 367 1114 387
rect 1118 367 1119 387
rect 504 320 505 340
rect 509 320 510 340
rect 679 320 680 340
rect 684 320 685 340
rect 854 320 855 340
rect 859 320 860 340
rect 1029 320 1030 340
rect 1034 320 1035 340
rect 2484 318 2485 338
rect 2489 318 2490 338
rect 2563 309 2564 329
rect 2568 309 2569 329
rect 2662 318 2663 338
rect 2667 318 2668 338
rect 2741 309 2742 329
rect 2746 309 2747 329
rect 2817 318 2818 338
rect 2822 318 2823 338
rect 2896 309 2897 329
rect 2901 309 2902 329
rect 2973 318 2974 338
rect 2978 318 2979 338
rect 3052 309 3053 329
rect 3057 309 3058 329
rect 2368 282 2369 302
rect 2373 282 2374 302
rect 658 187 659 207
rect 663 187 664 207
rect 742 194 743 214
rect 747 194 748 214
rect 828 187 829 207
rect 833 187 834 207
rect 912 194 913 214
rect 917 194 918 214
rect 1202 200 1203 220
rect 1207 200 1208 220
rect 1286 207 1287 227
rect 1291 207 1292 227
rect 1377 200 1378 220
rect 1382 200 1383 220
rect 1461 207 1462 227
rect 1466 207 1467 227
rect 1552 200 1553 220
rect 1557 200 1558 220
rect 1636 207 1637 227
rect 1641 207 1642 227
rect 1727 200 1728 220
rect 1732 200 1733 220
rect 1811 207 1812 227
rect 1816 207 1817 227
rect 2564 224 2565 244
rect 2569 224 2570 244
rect 2742 224 2743 244
rect 2747 224 2748 244
rect 2897 224 2898 244
rect 2902 224 2903 244
rect 3053 224 3054 244
rect 3058 224 3059 244
rect 573 147 574 167
rect 578 147 579 167
rect 658 147 659 167
rect 663 147 664 167
rect 828 147 829 167
rect 833 147 834 167
rect 1202 160 1203 180
rect 1207 160 1208 180
rect 1377 160 1378 180
rect 1382 160 1383 180
rect 1552 160 1553 180
rect 1557 160 1558 180
rect 1727 160 1728 180
rect 1732 160 1733 180
rect 2307 89 2308 109
rect 2312 89 2313 109
rect 2391 96 2392 116
rect 2396 96 2397 116
rect 2489 89 2490 109
rect 2494 89 2495 109
rect 2573 96 2574 116
rect 2578 96 2579 116
rect 2829 89 2830 109
rect 2834 89 2835 109
rect 2913 96 2914 116
rect 2918 96 2919 116
rect 3011 89 3012 109
rect 3016 89 3017 109
rect 3095 96 3096 116
rect 3100 96 3101 116
rect 658 49 659 69
rect 663 49 664 69
rect 742 56 743 76
rect 747 56 748 76
rect 828 49 829 69
rect 833 49 834 69
rect 912 56 913 76
rect 917 56 918 76
rect 1202 49 1203 69
rect 1207 49 1208 69
rect 1286 56 1287 76
rect 1291 56 1292 76
rect 1377 49 1378 69
rect 1382 49 1383 69
rect 1461 56 1462 76
rect 1466 56 1467 76
rect 1552 49 1553 69
rect 1557 49 1558 69
rect 1636 56 1637 76
rect 1641 56 1642 76
rect 1727 49 1728 69
rect 1732 49 1733 69
rect 1811 56 1812 76
rect 1816 56 1817 76
rect 2307 49 2308 69
rect 2312 49 2313 69
rect 2489 49 2490 69
rect 2494 49 2495 69
rect 2645 53 2646 73
rect 2650 53 2651 73
rect 2696 53 2697 73
rect 2701 53 2702 73
rect 2743 56 2744 76
rect 2748 56 2749 76
rect 2829 49 2830 69
rect 2834 49 2835 69
rect 3011 49 3012 69
rect 3016 49 3017 69
rect 3167 53 3168 73
rect 3172 53 3173 73
rect 3218 53 3219 73
rect 3223 53 3224 73
rect 3265 56 3266 76
rect 3270 56 3271 76
rect 573 9 574 29
rect 578 9 579 29
rect 658 9 659 29
rect 663 9 664 29
rect 828 9 829 29
rect 833 9 834 29
rect 1012 13 1013 33
rect 1017 13 1018 33
rect 1063 13 1064 33
rect 1068 13 1069 33
rect 1110 16 1111 36
rect 1115 16 1116 36
rect 1202 9 1203 29
rect 1207 9 1208 29
rect 1377 9 1378 29
rect 1382 9 1383 29
rect 1552 9 1553 29
rect 1557 9 1558 29
rect 1727 9 1728 29
rect 1732 9 1733 29
rect 2339 -33 2340 -13
rect 2344 -33 2345 -13
rect 2418 -42 2419 -22
rect 2423 -42 2424 -22
rect 2650 -30 2651 -10
rect 2655 -30 2656 -10
rect 2729 -39 2730 -19
rect 2734 -39 2735 -19
rect 2861 -33 2862 -13
rect 2866 -33 2867 -13
rect 2940 -42 2941 -22
rect 2945 -42 2946 -22
rect 3172 -30 3173 -10
rect 3177 -30 3178 -10
rect 3251 -39 3252 -19
rect 3256 -39 3257 -19
rect 2339 -115 2340 -95
rect 2344 -115 2345 -95
rect 2419 -127 2420 -107
rect 2424 -127 2425 -107
rect 2650 -112 2651 -92
rect 2655 -112 2656 -92
rect 2730 -124 2731 -104
rect 2735 -124 2736 -104
rect 2861 -115 2862 -95
rect 2866 -115 2867 -95
rect 2941 -127 2942 -107
rect 2946 -127 2947 -107
rect 3172 -112 3173 -92
rect 3177 -112 3178 -92
rect 3252 -124 3253 -104
rect 3257 -124 3258 -104
rect 547 -197 548 -177
rect 552 -197 553 -177
rect 631 -190 632 -170
rect 636 -190 637 -170
rect 722 -197 723 -177
rect 727 -197 728 -177
rect 806 -190 807 -170
rect 811 -190 812 -170
rect 897 -197 898 -177
rect 902 -197 903 -177
rect 981 -190 982 -170
rect 986 -190 987 -170
rect 1072 -197 1073 -177
rect 1077 -197 1078 -177
rect 1156 -190 1157 -170
rect 1161 -190 1162 -170
rect 547 -237 548 -217
rect 552 -237 553 -217
rect 722 -237 723 -217
rect 727 -237 728 -217
rect 897 -237 898 -217
rect 902 -237 903 -217
rect 1072 -237 1073 -217
rect 1077 -237 1078 -217
rect 2307 -297 2308 -277
rect 2312 -297 2313 -277
rect 2391 -290 2392 -270
rect 2396 -290 2397 -270
rect 2489 -297 2490 -277
rect 2494 -297 2495 -277
rect 2573 -290 2574 -270
rect 2578 -290 2579 -270
rect 2829 -297 2830 -277
rect 2834 -297 2835 -277
rect 2913 -290 2914 -270
rect 2918 -290 2919 -270
rect 3011 -297 3012 -277
rect 3016 -297 3017 -277
rect 3095 -290 3096 -270
rect 3100 -290 3101 -270
rect 547 -348 548 -328
rect 552 -348 553 -328
rect 631 -341 632 -321
rect 636 -341 637 -321
rect 722 -348 723 -328
rect 727 -348 728 -328
rect 806 -341 807 -321
rect 811 -341 812 -321
rect 897 -348 898 -328
rect 902 -348 903 -328
rect 981 -341 982 -321
rect 986 -341 987 -321
rect 1072 -348 1073 -328
rect 1077 -348 1078 -328
rect 1156 -341 1157 -321
rect 1161 -341 1162 -321
rect 2307 -337 2308 -317
rect 2312 -337 2313 -317
rect 2489 -337 2490 -317
rect 2494 -337 2495 -317
rect 2645 -333 2646 -313
rect 2650 -333 2651 -313
rect 2696 -333 2697 -313
rect 2701 -333 2702 -313
rect 2743 -330 2744 -310
rect 2748 -330 2749 -310
rect 2829 -337 2830 -317
rect 2834 -337 2835 -317
rect 3011 -337 3012 -317
rect 3016 -337 3017 -317
rect 3167 -333 3168 -313
rect 3172 -333 3173 -313
rect 3218 -333 3219 -313
rect 3223 -333 3224 -313
rect 3265 -330 3266 -310
rect 3270 -330 3271 -310
rect 547 -388 548 -368
rect 552 -388 553 -368
rect 722 -388 723 -368
rect 727 -388 728 -368
rect 897 -388 898 -368
rect 902 -388 903 -368
rect 1072 -388 1073 -368
rect 1077 -388 1078 -368
rect 2339 -419 2340 -399
rect 2344 -419 2345 -399
rect 2418 -428 2419 -408
rect 2423 -428 2424 -408
rect 2650 -416 2651 -396
rect 2655 -416 2656 -396
rect 2729 -425 2730 -405
rect 2734 -425 2735 -405
rect 2861 -419 2862 -399
rect 2866 -419 2867 -399
rect 2940 -428 2941 -408
rect 2945 -428 2946 -408
rect 3172 -416 3173 -396
rect 3177 -416 3178 -396
rect 3251 -425 3252 -405
rect 3256 -425 3257 -405
rect 643 -507 644 -487
rect 648 -507 649 -487
rect 722 -516 723 -496
rect 727 -516 728 -496
rect 784 -507 785 -487
rect 789 -507 790 -487
rect 863 -516 864 -496
rect 868 -516 869 -496
rect 955 -523 956 -503
rect 960 -523 961 -503
rect 1148 -516 1149 -496
rect 1153 -516 1154 -496
rect 2339 -501 2340 -481
rect 2344 -501 2345 -481
rect 2419 -513 2420 -493
rect 2424 -513 2425 -493
rect 2650 -498 2651 -478
rect 2655 -498 2656 -478
rect 2730 -510 2731 -490
rect 2735 -510 2736 -490
rect 2861 -501 2862 -481
rect 2866 -501 2867 -481
rect 2941 -513 2942 -493
rect 2946 -513 2947 -493
rect 3172 -498 3173 -478
rect 3177 -498 3178 -478
rect 3252 -510 3253 -490
rect 3257 -510 3258 -490
rect 955 -563 956 -543
rect 960 -563 961 -543
rect 643 -589 644 -569
rect 648 -589 649 -569
rect 723 -601 724 -581
rect 728 -601 729 -581
rect 784 -589 785 -569
rect 789 -589 790 -569
rect 864 -601 865 -581
rect 869 -601 870 -581
rect 955 -603 956 -583
rect 960 -603 961 -583
rect 1272 -588 1273 -568
rect 1277 -588 1278 -568
rect 955 -642 956 -622
rect 960 -642 961 -622
rect 1272 -628 1273 -608
rect 1277 -628 1278 -608
rect 1272 -668 1273 -648
rect 1277 -668 1278 -648
rect 1634 -659 1635 -639
rect 1639 -659 1640 -639
rect 1718 -652 1719 -632
rect 1723 -652 1724 -632
rect 1804 -659 1805 -639
rect 1809 -659 1810 -639
rect 1888 -652 1889 -632
rect 1893 -652 1894 -632
rect 1974 -659 1975 -639
rect 1979 -659 1980 -639
rect 2058 -652 2059 -632
rect 2063 -652 2064 -632
rect 2144 -659 2145 -639
rect 2149 -659 2150 -639
rect 2228 -652 2229 -632
rect 2233 -652 2234 -632
rect 643 -688 644 -668
rect 648 -688 649 -668
rect 722 -697 723 -677
rect 727 -697 728 -677
rect 784 -688 785 -668
rect 789 -688 790 -668
rect 863 -697 864 -677
rect 868 -697 869 -677
rect 1272 -707 1273 -687
rect 1277 -707 1278 -687
rect 1634 -699 1635 -679
rect 1639 -699 1640 -679
rect 1804 -699 1805 -679
rect 1809 -699 1810 -679
rect 1974 -699 1975 -679
rect 1979 -699 1980 -679
rect 2144 -699 2145 -679
rect 2149 -699 2150 -679
rect 985 -740 986 -720
rect 990 -740 991 -720
rect 1272 -746 1273 -726
rect 1277 -746 1278 -726
rect 643 -770 644 -750
rect 648 -770 649 -750
rect 723 -782 724 -762
rect 728 -782 729 -762
rect 784 -770 785 -750
rect 789 -770 790 -750
rect 864 -782 865 -762
rect 869 -782 870 -762
rect 985 -780 986 -760
rect 990 -780 991 -760
rect 1102 -780 1103 -760
rect 1107 -780 1108 -760
rect 1153 -780 1154 -760
rect 1158 -780 1159 -760
rect 670 -885 671 -865
rect 675 -885 676 -865
rect 878 -884 879 -864
rect 883 -884 884 -864
rect 1170 -884 1171 -864
rect 1175 -884 1176 -864
rect 670 -925 671 -905
rect 675 -925 676 -905
rect 878 -924 879 -904
rect 883 -924 884 -904
rect 1170 -924 1171 -904
rect 1175 -924 1176 -904
rect 670 -965 671 -945
rect 675 -965 676 -945
rect 878 -964 879 -944
rect 883 -964 884 -944
rect 1170 -964 1171 -944
rect 1175 -964 1176 -944
rect 1452 -962 1453 -942
rect 1457 -962 1458 -942
rect 1536 -955 1537 -935
rect 1541 -955 1542 -935
rect 878 -1003 879 -983
rect 883 -1003 884 -983
rect 1170 -1003 1171 -983
rect 1175 -1003 1176 -983
rect 1452 -1002 1453 -982
rect 1457 -1002 1458 -982
<< pdiffusion >>
rect 478 563 479 583
rect 481 563 482 583
rect 534 563 535 583
rect 537 563 538 583
rect 589 554 590 574
rect 592 554 593 574
rect 653 563 654 583
rect 656 563 657 583
rect 709 563 710 583
rect 712 563 713 583
rect 764 554 765 574
rect 767 554 768 574
rect 828 563 829 583
rect 831 563 832 583
rect 884 563 885 583
rect 887 563 888 583
rect 939 554 940 574
rect 942 554 943 574
rect 1003 563 1004 583
rect 1006 563 1007 583
rect 1059 563 1060 583
rect 1062 563 1063 583
rect 1114 554 1115 574
rect 1117 554 1118 574
rect 1181 563 1182 583
rect 1184 563 1185 583
rect 1237 563 1238 583
rect 1240 563 1241 583
rect 1292 554 1293 574
rect 1295 554 1296 574
rect 1351 563 1352 583
rect 1354 563 1355 583
rect 1407 563 1408 583
rect 1410 563 1411 583
rect 1462 554 1463 574
rect 1465 554 1466 574
rect 1521 563 1522 583
rect 1524 563 1525 583
rect 1577 563 1578 583
rect 1580 563 1581 583
rect 1632 554 1633 574
rect 1635 554 1636 574
rect 1691 563 1692 583
rect 1694 563 1695 583
rect 1747 563 1748 583
rect 1750 563 1751 583
rect 1802 554 1803 574
rect 1805 554 1806 574
rect 478 412 479 432
rect 481 412 482 432
rect 534 412 535 432
rect 537 412 538 432
rect 589 403 590 423
rect 592 403 593 423
rect 653 412 654 432
rect 656 412 657 432
rect 709 412 710 432
rect 712 412 713 432
rect 764 403 765 423
rect 767 403 768 423
rect 828 412 829 432
rect 831 412 832 432
rect 884 412 885 432
rect 887 412 888 432
rect 939 403 940 423
rect 942 403 943 423
rect 1003 412 1004 432
rect 1006 412 1007 432
rect 1059 412 1060 432
rect 1062 412 1063 432
rect 1114 403 1115 423
rect 1117 403 1118 423
rect 2485 354 2486 374
rect 2488 354 2489 374
rect 2548 354 2549 374
rect 2551 354 2552 374
rect 2663 354 2664 374
rect 2666 354 2667 374
rect 2726 354 2727 374
rect 2729 354 2730 374
rect 2818 354 2819 374
rect 2821 354 2822 374
rect 2881 354 2882 374
rect 2884 354 2885 374
rect 2974 354 2975 374
rect 2977 354 2978 374
rect 3037 354 3038 374
rect 3040 354 3041 374
rect 2369 318 2370 338
rect 2372 318 2373 338
rect 632 239 633 259
rect 635 239 636 259
rect 688 239 689 259
rect 691 239 692 259
rect 743 230 744 250
rect 746 230 747 250
rect 802 239 803 259
rect 805 239 806 259
rect 858 239 859 259
rect 861 239 862 259
rect 1176 252 1177 272
rect 1179 252 1180 272
rect 1232 252 1233 272
rect 1235 252 1236 272
rect 913 230 914 250
rect 916 230 917 250
rect 1287 243 1288 263
rect 1290 243 1291 263
rect 1351 252 1352 272
rect 1354 252 1355 272
rect 1407 252 1408 272
rect 1410 252 1411 272
rect 1462 243 1463 263
rect 1465 243 1466 263
rect 1526 252 1527 272
rect 1529 252 1530 272
rect 1582 252 1583 272
rect 1585 252 1586 272
rect 1637 243 1638 263
rect 1640 243 1641 263
rect 1701 252 1702 272
rect 1704 252 1705 272
rect 1757 252 1758 272
rect 1760 252 1761 272
rect 2549 269 2550 289
rect 2552 269 2553 289
rect 2727 269 2728 289
rect 2730 269 2731 289
rect 2882 269 2883 289
rect 2885 269 2886 289
rect 3038 269 3039 289
rect 3041 269 3042 289
rect 1812 243 1813 263
rect 1815 243 1816 263
rect 574 183 575 203
rect 577 183 578 203
rect 2281 141 2282 161
rect 2284 141 2285 161
rect 2337 141 2338 161
rect 2340 141 2341 161
rect 2392 132 2393 152
rect 2395 132 2396 152
rect 2463 141 2464 161
rect 2466 141 2467 161
rect 2519 141 2520 161
rect 2522 141 2523 161
rect 2574 132 2575 152
rect 2577 132 2578 152
rect 2656 145 2657 165
rect 2659 145 2660 165
rect 2803 141 2804 161
rect 2806 141 2807 161
rect 2859 141 2860 161
rect 2862 141 2863 161
rect 2914 132 2915 152
rect 2917 132 2918 152
rect 2985 141 2986 161
rect 2988 141 2989 161
rect 3041 141 3042 161
rect 3044 141 3045 161
rect 3096 132 3097 152
rect 3099 132 3100 152
rect 3178 145 3179 165
rect 3181 145 3182 165
rect 632 101 633 121
rect 635 101 636 121
rect 688 101 689 121
rect 691 101 692 121
rect 743 92 744 112
rect 746 92 747 112
rect 802 101 803 121
rect 805 101 806 121
rect 858 101 859 121
rect 861 101 862 121
rect 913 92 914 112
rect 916 92 917 112
rect 1023 105 1024 125
rect 1026 105 1027 125
rect 1176 101 1177 121
rect 1179 101 1180 121
rect 1232 101 1233 121
rect 1235 101 1236 121
rect 1287 92 1288 112
rect 1290 92 1291 112
rect 1351 101 1352 121
rect 1354 101 1355 121
rect 1407 101 1408 121
rect 1410 101 1411 121
rect 1462 92 1463 112
rect 1465 92 1466 112
rect 1526 101 1527 121
rect 1529 101 1530 121
rect 1582 101 1583 121
rect 1585 101 1586 121
rect 1637 92 1638 112
rect 1640 92 1641 112
rect 1701 101 1702 121
rect 1704 101 1705 121
rect 1757 101 1758 121
rect 1760 101 1761 121
rect 1812 92 1813 112
rect 1815 92 1816 112
rect 2656 99 2657 119
rect 2659 99 2660 119
rect 2744 92 2745 112
rect 2747 92 2748 112
rect 3178 99 3179 119
rect 3181 99 3182 119
rect 3266 92 3267 112
rect 3269 92 3270 112
rect 574 45 575 65
rect 577 45 578 65
rect 1023 59 1024 79
rect 1026 59 1027 79
rect 1111 52 1112 72
rect 1114 52 1115 72
rect 2340 3 2341 23
rect 2343 3 2344 23
rect 2403 3 2404 23
rect 2406 3 2407 23
rect 2651 6 2652 26
rect 2654 6 2655 26
rect 2714 6 2715 26
rect 2717 6 2718 26
rect 2862 3 2863 23
rect 2865 3 2866 23
rect 2925 3 2926 23
rect 2928 3 2929 23
rect 3173 6 3174 26
rect 3176 6 3177 26
rect 3236 6 3237 26
rect 3239 6 3240 26
rect 2340 -79 2341 -59
rect 2343 -79 2344 -59
rect 2404 -82 2405 -62
rect 2407 -82 2408 -62
rect 2651 -76 2652 -56
rect 2654 -76 2655 -56
rect 2715 -79 2716 -59
rect 2718 -79 2719 -59
rect 2862 -79 2863 -59
rect 2865 -79 2866 -59
rect 2926 -82 2927 -62
rect 2929 -82 2930 -62
rect 3173 -76 3174 -56
rect 3176 -76 3177 -56
rect 3237 -79 3238 -59
rect 3240 -79 3241 -59
rect 521 -145 522 -125
rect 524 -145 525 -125
rect 577 -145 578 -125
rect 580 -145 581 -125
rect 632 -154 633 -134
rect 635 -154 636 -134
rect 696 -145 697 -125
rect 699 -145 700 -125
rect 752 -145 753 -125
rect 755 -145 756 -125
rect 807 -154 808 -134
rect 810 -154 811 -134
rect 871 -145 872 -125
rect 874 -145 875 -125
rect 927 -145 928 -125
rect 930 -145 931 -125
rect 982 -154 983 -134
rect 985 -154 986 -134
rect 1046 -145 1047 -125
rect 1049 -145 1050 -125
rect 1102 -145 1103 -125
rect 1105 -145 1106 -125
rect 1157 -154 1158 -134
rect 1160 -154 1161 -134
rect 2281 -245 2282 -225
rect 2284 -245 2285 -225
rect 2337 -245 2338 -225
rect 2340 -245 2341 -225
rect 2392 -254 2393 -234
rect 2395 -254 2396 -234
rect 2463 -245 2464 -225
rect 2466 -245 2467 -225
rect 2519 -245 2520 -225
rect 2522 -245 2523 -225
rect 2574 -254 2575 -234
rect 2577 -254 2578 -234
rect 2656 -241 2657 -221
rect 2659 -241 2660 -221
rect 2803 -245 2804 -225
rect 2806 -245 2807 -225
rect 2859 -245 2860 -225
rect 2862 -245 2863 -225
rect 2914 -254 2915 -234
rect 2917 -254 2918 -234
rect 2985 -245 2986 -225
rect 2988 -245 2989 -225
rect 3041 -245 3042 -225
rect 3044 -245 3045 -225
rect 3096 -254 3097 -234
rect 3099 -254 3100 -234
rect 3178 -241 3179 -221
rect 3181 -241 3182 -221
rect 521 -296 522 -276
rect 524 -296 525 -276
rect 577 -296 578 -276
rect 580 -296 581 -276
rect 632 -305 633 -285
rect 635 -305 636 -285
rect 696 -296 697 -276
rect 699 -296 700 -276
rect 752 -296 753 -276
rect 755 -296 756 -276
rect 807 -305 808 -285
rect 810 -305 811 -285
rect 871 -296 872 -276
rect 874 -296 875 -276
rect 927 -296 928 -276
rect 930 -296 931 -276
rect 982 -305 983 -285
rect 985 -305 986 -285
rect 1046 -296 1047 -276
rect 1049 -296 1050 -276
rect 1102 -296 1103 -276
rect 1105 -296 1106 -276
rect 1157 -305 1158 -285
rect 1160 -305 1161 -285
rect 2656 -287 2657 -267
rect 2659 -287 2660 -267
rect 2744 -294 2745 -274
rect 2747 -294 2748 -274
rect 3178 -287 3179 -267
rect 3181 -287 3182 -267
rect 3266 -294 3267 -274
rect 3269 -294 3270 -274
rect 2340 -383 2341 -363
rect 2343 -383 2344 -363
rect 2403 -383 2404 -363
rect 2406 -383 2407 -363
rect 2651 -380 2652 -360
rect 2654 -380 2655 -360
rect 2714 -380 2715 -360
rect 2717 -380 2718 -360
rect 2862 -383 2863 -363
rect 2865 -383 2866 -363
rect 2925 -383 2926 -363
rect 2928 -383 2929 -363
rect 3173 -380 3174 -360
rect 3176 -380 3177 -360
rect 3236 -380 3237 -360
rect 3239 -380 3240 -360
rect 644 -471 645 -451
rect 647 -471 648 -451
rect 707 -471 708 -451
rect 710 -471 711 -451
rect 785 -471 786 -451
rect 788 -471 789 -451
rect 848 -471 849 -451
rect 851 -471 852 -451
rect 929 -471 930 -451
rect 932 -471 933 -451
rect 985 -471 986 -451
rect 988 -471 989 -451
rect 1041 -471 1042 -451
rect 1044 -471 1045 -451
rect 1097 -471 1098 -451
rect 1100 -471 1101 -451
rect 1149 -480 1150 -460
rect 1152 -480 1153 -460
rect 2340 -465 2341 -445
rect 2343 -465 2344 -445
rect 2404 -468 2405 -448
rect 2407 -468 2408 -448
rect 2651 -462 2652 -442
rect 2654 -462 2655 -442
rect 2715 -465 2716 -445
rect 2718 -465 2719 -445
rect 2862 -465 2863 -445
rect 2865 -465 2866 -445
rect 2926 -468 2927 -448
rect 2929 -468 2930 -448
rect 3173 -462 3174 -442
rect 3176 -462 3177 -442
rect 3237 -465 3238 -445
rect 3240 -465 3241 -445
rect 644 -553 645 -533
rect 647 -553 648 -533
rect 708 -556 709 -536
rect 711 -556 712 -536
rect 785 -553 786 -533
rect 788 -553 789 -533
rect 1246 -536 1247 -516
rect 1249 -536 1250 -516
rect 1302 -536 1303 -516
rect 1305 -536 1306 -516
rect 1358 -536 1359 -516
rect 1361 -536 1362 -516
rect 1414 -536 1415 -516
rect 1417 -536 1418 -516
rect 1469 -536 1470 -516
rect 1472 -536 1473 -516
rect 849 -556 850 -536
rect 852 -556 853 -536
rect 1608 -607 1609 -587
rect 1611 -607 1612 -587
rect 1664 -607 1665 -587
rect 1667 -607 1668 -587
rect 644 -652 645 -632
rect 647 -652 648 -632
rect 707 -652 708 -632
rect 710 -652 711 -632
rect 785 -652 786 -632
rect 788 -652 789 -632
rect 848 -652 849 -632
rect 851 -652 852 -632
rect 1719 -616 1720 -596
rect 1722 -616 1723 -596
rect 1778 -607 1779 -587
rect 1781 -607 1782 -587
rect 1834 -607 1835 -587
rect 1837 -607 1838 -587
rect 1889 -616 1890 -596
rect 1892 -616 1893 -596
rect 1948 -607 1949 -587
rect 1951 -607 1952 -587
rect 2004 -607 2005 -587
rect 2007 -607 2008 -587
rect 2059 -616 2060 -596
rect 2062 -616 2063 -596
rect 2118 -607 2119 -587
rect 2121 -607 2122 -587
rect 2174 -607 2175 -587
rect 2177 -607 2178 -587
rect 2229 -616 2230 -596
rect 2232 -616 2233 -596
rect 959 -688 960 -668
rect 962 -688 963 -668
rect 1015 -688 1016 -668
rect 1018 -688 1019 -668
rect 1113 -688 1114 -668
rect 1116 -688 1117 -668
rect 644 -734 645 -714
rect 647 -734 648 -714
rect 708 -737 709 -717
rect 711 -737 712 -717
rect 785 -734 786 -714
rect 788 -734 789 -714
rect 849 -737 850 -717
rect 852 -737 853 -717
rect 1113 -734 1114 -714
rect 1116 -734 1117 -714
rect 644 -833 645 -813
rect 647 -833 648 -813
rect 700 -833 701 -813
rect 703 -833 704 -813
rect 756 -833 757 -813
rect 759 -833 760 -813
rect 852 -832 853 -812
rect 855 -832 856 -812
rect 908 -832 909 -812
rect 911 -832 912 -812
rect 964 -832 965 -812
rect 967 -832 968 -812
rect 1020 -832 1021 -812
rect 1023 -832 1024 -812
rect 1144 -832 1145 -812
rect 1147 -832 1148 -812
rect 1200 -832 1201 -812
rect 1203 -832 1204 -812
rect 1256 -832 1257 -812
rect 1259 -832 1260 -812
rect 1312 -832 1313 -812
rect 1315 -832 1316 -812
rect 1426 -910 1427 -890
rect 1429 -910 1430 -890
rect 1482 -910 1483 -890
rect 1485 -910 1486 -890
rect 1537 -919 1538 -899
rect 1540 -919 1541 -899
<< ndcontact >>
rect 494 511 504 531
rect 510 511 520 531
rect 578 518 588 538
rect 594 518 604 538
rect 669 511 679 531
rect 685 511 695 531
rect 753 518 763 538
rect 769 518 779 538
rect 844 511 854 531
rect 860 511 870 531
rect 928 518 938 538
rect 944 518 954 538
rect 1019 511 1029 531
rect 1035 511 1045 531
rect 1103 518 1113 538
rect 1119 518 1129 538
rect 1197 511 1207 531
rect 1213 511 1223 531
rect 1281 518 1291 538
rect 1297 518 1307 538
rect 1367 511 1377 531
rect 1383 511 1393 531
rect 1451 518 1461 538
rect 1467 518 1477 538
rect 1537 511 1547 531
rect 1553 511 1563 531
rect 1621 518 1631 538
rect 1637 518 1647 538
rect 1707 511 1717 531
rect 1723 511 1733 531
rect 1791 518 1801 538
rect 1807 518 1817 538
rect 494 471 504 491
rect 510 471 520 491
rect 669 471 679 491
rect 685 471 695 491
rect 844 471 854 491
rect 860 471 870 491
rect 1019 471 1029 491
rect 1035 471 1045 491
rect 1197 471 1207 491
rect 1213 471 1223 491
rect 1367 471 1377 491
rect 1383 471 1393 491
rect 1537 471 1547 491
rect 1553 471 1563 491
rect 1707 471 1717 491
rect 1723 471 1733 491
rect 494 360 504 380
rect 510 360 520 380
rect 578 367 588 387
rect 594 367 604 387
rect 669 360 679 380
rect 685 360 695 380
rect 753 367 763 387
rect 769 367 779 387
rect 844 360 854 380
rect 860 360 870 380
rect 928 367 938 387
rect 944 367 954 387
rect 1019 360 1029 380
rect 1035 360 1045 380
rect 1103 367 1113 387
rect 1119 367 1129 387
rect 494 320 504 340
rect 510 320 520 340
rect 669 320 679 340
rect 685 320 695 340
rect 844 320 854 340
rect 860 320 870 340
rect 1019 320 1029 340
rect 1035 320 1045 340
rect 2474 318 2484 338
rect 2490 318 2500 338
rect 2553 309 2563 329
rect 2569 309 2579 329
rect 2652 318 2662 338
rect 2668 318 2678 338
rect 2731 309 2741 329
rect 2747 309 2757 329
rect 2807 318 2817 338
rect 2823 318 2833 338
rect 2886 309 2896 329
rect 2902 309 2912 329
rect 2963 318 2973 338
rect 2979 318 2989 338
rect 3042 309 3052 329
rect 3058 309 3068 329
rect 2358 282 2368 302
rect 2374 282 2384 302
rect 648 187 658 207
rect 664 187 674 207
rect 732 194 742 214
rect 748 194 758 214
rect 818 187 828 207
rect 834 187 844 207
rect 902 194 912 214
rect 918 194 928 214
rect 1192 200 1202 220
rect 1208 200 1218 220
rect 1276 207 1286 227
rect 1292 207 1302 227
rect 1367 200 1377 220
rect 1383 200 1393 220
rect 1451 207 1461 227
rect 1467 207 1477 227
rect 1542 200 1552 220
rect 1558 200 1568 220
rect 1626 207 1636 227
rect 1642 207 1652 227
rect 1717 200 1727 220
rect 1733 200 1743 220
rect 1801 207 1811 227
rect 1817 207 1827 227
rect 2554 224 2564 244
rect 2570 224 2579 244
rect 2732 224 2742 244
rect 2748 224 2757 244
rect 2887 224 2897 244
rect 2903 224 2912 244
rect 3043 224 3053 244
rect 3059 224 3068 244
rect 563 147 573 167
rect 579 147 589 167
rect 648 147 658 167
rect 664 147 674 167
rect 818 147 828 167
rect 834 147 844 167
rect 1192 160 1202 180
rect 1208 160 1218 180
rect 1367 160 1377 180
rect 1383 160 1393 180
rect 1542 160 1552 180
rect 1558 160 1568 180
rect 1717 160 1727 180
rect 1733 160 1743 180
rect 2297 89 2307 109
rect 2313 89 2323 109
rect 2381 96 2391 116
rect 2397 96 2407 116
rect 2479 89 2489 109
rect 2495 89 2505 109
rect 2563 96 2573 116
rect 2579 96 2589 116
rect 2819 89 2829 109
rect 2835 89 2845 109
rect 2903 96 2913 116
rect 2919 96 2929 116
rect 3001 89 3011 109
rect 3017 89 3027 109
rect 3085 96 3095 116
rect 3101 96 3111 116
rect 648 49 658 69
rect 664 49 674 69
rect 732 56 742 76
rect 748 56 758 76
rect 818 49 828 69
rect 834 49 844 69
rect 902 56 912 76
rect 918 56 928 76
rect 1192 49 1202 69
rect 1208 49 1218 69
rect 1276 56 1286 76
rect 1292 56 1302 76
rect 1367 49 1377 69
rect 1383 49 1393 69
rect 1451 56 1461 76
rect 1467 56 1477 76
rect 1542 49 1552 69
rect 1558 49 1568 69
rect 1626 56 1636 76
rect 1642 56 1652 76
rect 1717 49 1727 69
rect 1733 49 1743 69
rect 1801 56 1811 76
rect 1817 56 1827 76
rect 2297 49 2307 69
rect 2313 49 2323 69
rect 2479 49 2489 69
rect 2495 49 2505 69
rect 2635 53 2645 73
rect 2651 53 2661 73
rect 2686 53 2696 73
rect 2702 53 2712 73
rect 2733 56 2743 76
rect 2749 56 2759 76
rect 2819 49 2829 69
rect 2835 49 2845 69
rect 3001 49 3011 69
rect 3017 49 3027 69
rect 3157 53 3167 73
rect 3173 53 3183 73
rect 3208 53 3218 73
rect 3224 53 3234 73
rect 3255 56 3265 76
rect 3271 56 3281 76
rect 563 9 573 29
rect 579 9 589 29
rect 648 9 658 29
rect 664 9 674 29
rect 818 9 828 29
rect 834 9 844 29
rect 1002 13 1012 33
rect 1018 13 1028 33
rect 1053 13 1063 33
rect 1069 13 1079 33
rect 1100 16 1110 36
rect 1116 16 1126 36
rect 1192 9 1202 29
rect 1208 9 1218 29
rect 1367 9 1377 29
rect 1383 9 1393 29
rect 1542 9 1552 29
rect 1558 9 1568 29
rect 1717 9 1727 29
rect 1733 9 1743 29
rect 2329 -33 2339 -13
rect 2345 -33 2355 -13
rect 2408 -42 2418 -22
rect 2424 -42 2434 -22
rect 2640 -30 2650 -10
rect 2656 -30 2666 -10
rect 2719 -39 2729 -19
rect 2735 -39 2745 -19
rect 2851 -33 2861 -13
rect 2867 -33 2877 -13
rect 2930 -42 2940 -22
rect 2946 -42 2956 -22
rect 3162 -30 3172 -10
rect 3178 -30 3188 -10
rect 3241 -39 3251 -19
rect 3257 -39 3267 -19
rect 2329 -115 2339 -95
rect 2345 -115 2355 -95
rect 2409 -127 2419 -107
rect 2425 -127 2434 -107
rect 2640 -112 2650 -92
rect 2656 -112 2666 -92
rect 2720 -124 2730 -104
rect 2736 -124 2745 -104
rect 2851 -115 2861 -95
rect 2867 -115 2877 -95
rect 2931 -127 2941 -107
rect 2947 -127 2956 -107
rect 3162 -112 3172 -92
rect 3178 -112 3188 -92
rect 3242 -124 3252 -104
rect 3258 -124 3267 -104
rect 537 -197 547 -177
rect 553 -197 563 -177
rect 621 -190 631 -170
rect 637 -190 647 -170
rect 712 -197 722 -177
rect 728 -197 738 -177
rect 796 -190 806 -170
rect 812 -190 822 -170
rect 887 -197 897 -177
rect 903 -197 913 -177
rect 971 -190 981 -170
rect 987 -190 997 -170
rect 1062 -197 1072 -177
rect 1078 -197 1088 -177
rect 1146 -190 1156 -170
rect 1162 -190 1172 -170
rect 537 -237 547 -217
rect 553 -237 563 -217
rect 712 -237 722 -217
rect 728 -237 738 -217
rect 887 -237 897 -217
rect 903 -237 913 -217
rect 1062 -237 1072 -217
rect 1078 -237 1088 -217
rect 2297 -297 2307 -277
rect 2313 -297 2323 -277
rect 2381 -290 2391 -270
rect 2397 -290 2407 -270
rect 2479 -297 2489 -277
rect 2495 -297 2505 -277
rect 2563 -290 2573 -270
rect 2579 -290 2589 -270
rect 2819 -297 2829 -277
rect 2835 -297 2845 -277
rect 2903 -290 2913 -270
rect 2919 -290 2929 -270
rect 3001 -297 3011 -277
rect 3017 -297 3027 -277
rect 3085 -290 3095 -270
rect 3101 -290 3111 -270
rect 537 -348 547 -328
rect 553 -348 563 -328
rect 621 -341 631 -321
rect 637 -341 647 -321
rect 712 -348 722 -328
rect 728 -348 738 -328
rect 796 -341 806 -321
rect 812 -341 822 -321
rect 887 -348 897 -328
rect 903 -348 913 -328
rect 971 -341 981 -321
rect 987 -341 997 -321
rect 1062 -348 1072 -328
rect 1078 -348 1088 -328
rect 1146 -341 1156 -321
rect 1162 -341 1172 -321
rect 2297 -337 2307 -317
rect 2313 -337 2323 -317
rect 2479 -337 2489 -317
rect 2495 -337 2505 -317
rect 2635 -333 2645 -313
rect 2651 -333 2661 -313
rect 2686 -333 2696 -313
rect 2702 -333 2712 -313
rect 2733 -330 2743 -310
rect 2749 -330 2759 -310
rect 2819 -337 2829 -317
rect 2835 -337 2845 -317
rect 3001 -337 3011 -317
rect 3017 -337 3027 -317
rect 3157 -333 3167 -313
rect 3173 -333 3183 -313
rect 3208 -333 3218 -313
rect 3224 -333 3234 -313
rect 3255 -330 3265 -310
rect 3271 -330 3281 -310
rect 537 -388 547 -368
rect 553 -388 563 -368
rect 712 -388 722 -368
rect 728 -388 738 -368
rect 887 -388 897 -368
rect 903 -388 913 -368
rect 1062 -388 1072 -368
rect 1078 -388 1088 -368
rect 2329 -419 2339 -399
rect 2345 -419 2355 -399
rect 2408 -428 2418 -408
rect 2424 -428 2434 -408
rect 2640 -416 2650 -396
rect 2656 -416 2666 -396
rect 2719 -425 2729 -405
rect 2735 -425 2745 -405
rect 2851 -419 2861 -399
rect 2867 -419 2877 -399
rect 2930 -428 2940 -408
rect 2946 -428 2956 -408
rect 3162 -416 3172 -396
rect 3178 -416 3188 -396
rect 3241 -425 3251 -405
rect 3257 -425 3267 -405
rect 633 -507 643 -487
rect 649 -507 659 -487
rect 712 -516 722 -496
rect 728 -516 738 -496
rect 774 -507 784 -487
rect 790 -507 800 -487
rect 853 -516 863 -496
rect 869 -516 879 -496
rect 945 -523 955 -503
rect 961 -523 971 -503
rect 1138 -516 1148 -496
rect 1154 -516 1164 -496
rect 2329 -501 2339 -481
rect 2345 -501 2355 -481
rect 2409 -513 2419 -493
rect 2425 -513 2434 -493
rect 2640 -498 2650 -478
rect 2656 -498 2666 -478
rect 2720 -510 2730 -490
rect 2736 -510 2745 -490
rect 2851 -501 2861 -481
rect 2867 -501 2877 -481
rect 2931 -513 2941 -493
rect 2947 -513 2956 -493
rect 3162 -498 3172 -478
rect 3178 -498 3188 -478
rect 3242 -510 3252 -490
rect 3258 -510 3267 -490
rect 945 -563 955 -543
rect 961 -563 971 -543
rect 633 -589 643 -569
rect 649 -589 659 -569
rect 713 -601 723 -581
rect 729 -601 738 -581
rect 774 -589 784 -569
rect 790 -589 800 -569
rect 854 -601 864 -581
rect 870 -601 879 -581
rect 945 -603 955 -583
rect 961 -603 971 -583
rect 1262 -588 1272 -568
rect 1278 -588 1288 -568
rect 945 -642 955 -622
rect 961 -642 971 -622
rect 1262 -628 1272 -608
rect 1278 -628 1288 -608
rect 1262 -668 1272 -648
rect 1278 -668 1288 -648
rect 1624 -659 1634 -639
rect 1640 -659 1650 -639
rect 1708 -652 1718 -632
rect 1724 -652 1734 -632
rect 1794 -659 1804 -639
rect 1810 -659 1820 -639
rect 1878 -652 1888 -632
rect 1894 -652 1904 -632
rect 1964 -659 1974 -639
rect 1980 -659 1990 -639
rect 2048 -652 2058 -632
rect 2064 -652 2074 -632
rect 2134 -659 2144 -639
rect 2150 -659 2160 -639
rect 2218 -652 2228 -632
rect 2234 -652 2244 -632
rect 633 -688 643 -668
rect 649 -688 659 -668
rect 712 -697 722 -677
rect 728 -697 738 -677
rect 774 -688 784 -668
rect 790 -688 800 -668
rect 853 -697 863 -677
rect 869 -697 879 -677
rect 1262 -707 1272 -687
rect 1278 -707 1288 -687
rect 1624 -699 1634 -679
rect 1640 -699 1650 -679
rect 1794 -699 1804 -679
rect 1810 -699 1820 -679
rect 1964 -699 1974 -679
rect 1980 -699 1990 -679
rect 2134 -699 2144 -679
rect 2150 -699 2160 -679
rect 975 -740 985 -720
rect 991 -740 1001 -720
rect 1262 -746 1272 -726
rect 1278 -746 1288 -726
rect 633 -770 643 -750
rect 649 -770 659 -750
rect 713 -782 723 -762
rect 729 -782 738 -762
rect 774 -770 784 -750
rect 790 -770 800 -750
rect 854 -782 864 -762
rect 870 -782 879 -762
rect 975 -780 985 -760
rect 991 -780 1001 -760
rect 1092 -780 1102 -760
rect 1108 -780 1118 -760
rect 1143 -780 1153 -760
rect 1159 -780 1169 -760
rect 660 -885 670 -865
rect 676 -885 686 -865
rect 868 -884 878 -864
rect 884 -884 894 -864
rect 1160 -884 1170 -864
rect 1176 -884 1186 -864
rect 660 -925 670 -905
rect 676 -925 686 -905
rect 868 -924 878 -904
rect 884 -924 894 -904
rect 1160 -924 1170 -904
rect 1176 -924 1186 -904
rect 660 -965 670 -945
rect 676 -965 686 -945
rect 868 -964 878 -944
rect 884 -964 894 -944
rect 1160 -964 1170 -944
rect 1176 -964 1186 -944
rect 1442 -962 1452 -942
rect 1458 -962 1468 -942
rect 1526 -955 1536 -935
rect 1542 -955 1552 -935
rect 868 -1003 878 -983
rect 884 -1003 894 -983
rect 1160 -1003 1170 -983
rect 1176 -1003 1186 -983
rect 1442 -1002 1452 -982
rect 1458 -1002 1468 -982
<< pdcontact >>
rect 468 563 478 583
rect 482 563 492 583
rect 524 563 534 583
rect 538 563 548 583
rect 579 554 589 574
rect 593 554 603 574
rect 643 563 653 583
rect 657 563 667 583
rect 699 563 709 583
rect 713 563 723 583
rect 754 554 764 574
rect 768 554 778 574
rect 818 563 828 583
rect 832 563 842 583
rect 874 563 884 583
rect 888 563 898 583
rect 929 554 939 574
rect 943 554 953 574
rect 993 563 1003 583
rect 1007 563 1017 583
rect 1049 563 1059 583
rect 1063 563 1073 583
rect 1104 554 1114 574
rect 1118 554 1128 574
rect 1171 563 1181 583
rect 1185 563 1195 583
rect 1227 563 1237 583
rect 1241 563 1251 583
rect 1282 554 1292 574
rect 1296 554 1306 574
rect 1341 563 1351 583
rect 1355 563 1365 583
rect 1397 563 1407 583
rect 1411 563 1421 583
rect 1452 554 1462 574
rect 1466 554 1476 574
rect 1511 563 1521 583
rect 1525 563 1535 583
rect 1567 563 1577 583
rect 1581 563 1591 583
rect 1622 554 1632 574
rect 1636 554 1646 574
rect 1681 563 1691 583
rect 1695 563 1705 583
rect 1737 563 1747 583
rect 1751 563 1761 583
rect 1792 554 1802 574
rect 1806 554 1816 574
rect 468 412 478 432
rect 482 412 492 432
rect 524 412 534 432
rect 538 412 548 432
rect 579 403 589 423
rect 593 403 603 423
rect 643 412 653 432
rect 657 412 667 432
rect 699 412 709 432
rect 713 412 723 432
rect 754 403 764 423
rect 768 403 778 423
rect 818 412 828 432
rect 832 412 842 432
rect 874 412 884 432
rect 888 412 898 432
rect 929 403 939 423
rect 943 403 953 423
rect 993 412 1003 432
rect 1007 412 1017 432
rect 1049 412 1059 432
rect 1063 412 1073 432
rect 1104 403 1114 423
rect 1118 403 1128 423
rect 2475 354 2485 374
rect 2489 354 2499 374
rect 2538 354 2548 374
rect 2552 354 2562 374
rect 2653 354 2663 374
rect 2667 354 2677 374
rect 2716 354 2726 374
rect 2730 354 2740 374
rect 2808 354 2818 374
rect 2822 354 2832 374
rect 2871 354 2881 374
rect 2885 354 2895 374
rect 2964 354 2974 374
rect 2978 354 2988 374
rect 3027 354 3037 374
rect 3041 354 3051 374
rect 2359 318 2369 338
rect 2373 318 2383 338
rect 622 239 632 259
rect 636 239 646 259
rect 678 239 688 259
rect 692 239 702 259
rect 733 230 743 250
rect 747 230 757 250
rect 792 239 802 259
rect 806 239 816 259
rect 848 239 858 259
rect 862 239 872 259
rect 1166 252 1176 272
rect 1180 252 1190 272
rect 1222 252 1232 272
rect 1236 252 1246 272
rect 903 230 913 250
rect 917 230 927 250
rect 1277 243 1287 263
rect 1291 243 1301 263
rect 1341 252 1351 272
rect 1355 252 1365 272
rect 1397 252 1407 272
rect 1411 252 1421 272
rect 1452 243 1462 263
rect 1466 243 1476 263
rect 1516 252 1526 272
rect 1530 252 1540 272
rect 1572 252 1582 272
rect 1586 252 1596 272
rect 1627 243 1637 263
rect 1641 243 1651 263
rect 1691 252 1701 272
rect 1705 252 1715 272
rect 1747 252 1757 272
rect 1761 252 1771 272
rect 2539 269 2549 289
rect 2553 269 2563 289
rect 2717 269 2727 289
rect 2731 269 2741 289
rect 2872 269 2882 289
rect 2886 269 2896 289
rect 3028 269 3038 289
rect 3042 269 3052 289
rect 1802 243 1812 263
rect 1816 243 1826 263
rect 564 183 574 203
rect 578 183 588 203
rect 2271 141 2281 161
rect 2285 141 2295 161
rect 2327 141 2337 161
rect 2341 141 2351 161
rect 2382 132 2392 152
rect 2396 132 2406 152
rect 2453 141 2463 161
rect 2467 141 2477 161
rect 2509 141 2519 161
rect 2523 141 2533 161
rect 2564 132 2574 152
rect 2578 132 2588 152
rect 2646 145 2656 165
rect 2660 145 2670 165
rect 2793 141 2803 161
rect 2807 141 2817 161
rect 2849 141 2859 161
rect 2863 141 2873 161
rect 2904 132 2914 152
rect 2918 132 2928 152
rect 2975 141 2985 161
rect 2989 141 2999 161
rect 3031 141 3041 161
rect 3045 141 3055 161
rect 3086 132 3096 152
rect 3100 132 3110 152
rect 3168 145 3178 165
rect 3182 145 3192 165
rect 622 101 632 121
rect 636 101 646 121
rect 678 101 688 121
rect 692 101 702 121
rect 733 92 743 112
rect 747 92 757 112
rect 792 101 802 121
rect 806 101 816 121
rect 848 101 858 121
rect 862 101 872 121
rect 903 92 913 112
rect 917 92 927 112
rect 1013 105 1023 125
rect 1027 105 1037 125
rect 1166 101 1176 121
rect 1180 101 1190 121
rect 1222 101 1232 121
rect 1236 101 1246 121
rect 1277 92 1287 112
rect 1291 92 1301 112
rect 1341 101 1351 121
rect 1355 101 1365 121
rect 1397 101 1407 121
rect 1411 101 1421 121
rect 1452 92 1462 112
rect 1466 92 1476 112
rect 1516 101 1526 121
rect 1530 101 1540 121
rect 1572 101 1582 121
rect 1586 101 1596 121
rect 1627 92 1637 112
rect 1641 92 1651 112
rect 1691 101 1701 121
rect 1705 101 1715 121
rect 1747 101 1757 121
rect 1761 101 1771 121
rect 1802 92 1812 112
rect 1816 92 1826 112
rect 2646 99 2656 119
rect 2660 99 2670 119
rect 2734 92 2744 112
rect 2748 92 2758 112
rect 3168 99 3178 119
rect 3182 99 3192 119
rect 3256 92 3266 112
rect 3270 92 3280 112
rect 564 45 574 65
rect 578 45 588 65
rect 1013 59 1023 79
rect 1027 59 1037 79
rect 1101 52 1111 72
rect 1115 52 1125 72
rect 2330 3 2340 23
rect 2344 3 2354 23
rect 2393 3 2403 23
rect 2407 3 2417 23
rect 2641 6 2651 26
rect 2655 6 2665 26
rect 2704 6 2714 26
rect 2718 6 2728 26
rect 2852 3 2862 23
rect 2866 3 2876 23
rect 2915 3 2925 23
rect 2929 3 2939 23
rect 3163 6 3173 26
rect 3177 6 3187 26
rect 3226 6 3236 26
rect 3240 6 3250 26
rect 2330 -79 2340 -59
rect 2344 -79 2354 -59
rect 2394 -82 2404 -62
rect 2408 -82 2418 -62
rect 2641 -76 2651 -56
rect 2655 -76 2665 -56
rect 2705 -79 2715 -59
rect 2719 -79 2729 -59
rect 2852 -79 2862 -59
rect 2866 -79 2876 -59
rect 2916 -82 2926 -62
rect 2930 -82 2940 -62
rect 3163 -76 3173 -56
rect 3177 -76 3187 -56
rect 3227 -79 3237 -59
rect 3241 -79 3251 -59
rect 511 -145 521 -125
rect 525 -145 535 -125
rect 567 -145 577 -125
rect 581 -145 591 -125
rect 622 -154 632 -134
rect 636 -154 646 -134
rect 686 -145 696 -125
rect 700 -145 710 -125
rect 742 -145 752 -125
rect 756 -145 766 -125
rect 797 -154 807 -134
rect 811 -154 821 -134
rect 861 -145 871 -125
rect 875 -145 885 -125
rect 917 -145 927 -125
rect 931 -145 941 -125
rect 972 -154 982 -134
rect 986 -154 996 -134
rect 1036 -145 1046 -125
rect 1050 -145 1060 -125
rect 1092 -145 1102 -125
rect 1106 -145 1116 -125
rect 1147 -154 1157 -134
rect 1161 -154 1171 -134
rect 2271 -245 2281 -225
rect 2285 -245 2295 -225
rect 2327 -245 2337 -225
rect 2341 -245 2351 -225
rect 2382 -254 2392 -234
rect 2396 -254 2406 -234
rect 2453 -245 2463 -225
rect 2467 -245 2477 -225
rect 2509 -245 2519 -225
rect 2523 -245 2533 -225
rect 2564 -254 2574 -234
rect 2578 -254 2588 -234
rect 2646 -241 2656 -221
rect 2660 -241 2670 -221
rect 2793 -245 2803 -225
rect 2807 -245 2817 -225
rect 2849 -245 2859 -225
rect 2863 -245 2873 -225
rect 2904 -254 2914 -234
rect 2918 -254 2928 -234
rect 2975 -245 2985 -225
rect 2989 -245 2999 -225
rect 3031 -245 3041 -225
rect 3045 -245 3055 -225
rect 3086 -254 3096 -234
rect 3100 -254 3110 -234
rect 3168 -241 3178 -221
rect 3182 -241 3192 -221
rect 511 -296 521 -276
rect 525 -296 535 -276
rect 567 -296 577 -276
rect 581 -296 591 -276
rect 622 -305 632 -285
rect 636 -305 646 -285
rect 686 -296 696 -276
rect 700 -296 710 -276
rect 742 -296 752 -276
rect 756 -296 766 -276
rect 797 -305 807 -285
rect 811 -305 821 -285
rect 861 -296 871 -276
rect 875 -296 885 -276
rect 917 -296 927 -276
rect 931 -296 941 -276
rect 972 -305 982 -285
rect 986 -305 996 -285
rect 1036 -296 1046 -276
rect 1050 -296 1060 -276
rect 1092 -296 1102 -276
rect 1106 -296 1116 -276
rect 1147 -305 1157 -285
rect 1161 -305 1171 -285
rect 2646 -287 2656 -267
rect 2660 -287 2670 -267
rect 2734 -294 2744 -274
rect 2748 -294 2758 -274
rect 3168 -287 3178 -267
rect 3182 -287 3192 -267
rect 3256 -294 3266 -274
rect 3270 -294 3280 -274
rect 2330 -383 2340 -363
rect 2344 -383 2354 -363
rect 2393 -383 2403 -363
rect 2407 -383 2417 -363
rect 2641 -380 2651 -360
rect 2655 -380 2665 -360
rect 2704 -380 2714 -360
rect 2718 -380 2728 -360
rect 2852 -383 2862 -363
rect 2866 -383 2876 -363
rect 2915 -383 2925 -363
rect 2929 -383 2939 -363
rect 3163 -380 3173 -360
rect 3177 -380 3187 -360
rect 3226 -380 3236 -360
rect 3240 -380 3250 -360
rect 634 -471 644 -451
rect 648 -471 658 -451
rect 697 -471 707 -451
rect 711 -471 721 -451
rect 775 -471 785 -451
rect 789 -471 799 -451
rect 838 -471 848 -451
rect 852 -471 862 -451
rect 919 -471 929 -451
rect 933 -471 943 -451
rect 975 -471 985 -451
rect 989 -471 999 -451
rect 1031 -471 1041 -451
rect 1045 -471 1055 -451
rect 1087 -471 1097 -451
rect 1101 -471 1111 -451
rect 1139 -480 1149 -460
rect 1153 -480 1163 -460
rect 2330 -465 2340 -445
rect 2344 -465 2354 -445
rect 2394 -468 2404 -448
rect 2408 -468 2418 -448
rect 2641 -462 2651 -442
rect 2655 -462 2665 -442
rect 2705 -465 2715 -445
rect 2719 -465 2729 -445
rect 2852 -465 2862 -445
rect 2866 -465 2876 -445
rect 2916 -468 2926 -448
rect 2930 -468 2940 -448
rect 3163 -462 3173 -442
rect 3177 -462 3187 -442
rect 3227 -465 3237 -445
rect 3241 -465 3251 -445
rect 634 -553 644 -533
rect 648 -553 658 -533
rect 698 -556 708 -536
rect 712 -556 722 -536
rect 775 -553 785 -533
rect 789 -553 799 -533
rect 1236 -536 1246 -516
rect 1250 -536 1260 -516
rect 1292 -536 1302 -516
rect 1306 -536 1316 -516
rect 1348 -536 1358 -516
rect 1362 -536 1372 -516
rect 1404 -536 1414 -516
rect 1418 -536 1428 -516
rect 1459 -536 1469 -516
rect 1473 -536 1483 -516
rect 839 -556 849 -536
rect 853 -556 863 -536
rect 1598 -607 1608 -587
rect 1612 -607 1622 -587
rect 1654 -607 1664 -587
rect 1668 -607 1678 -587
rect 634 -652 644 -632
rect 648 -652 658 -632
rect 697 -652 707 -632
rect 711 -652 721 -632
rect 775 -652 785 -632
rect 789 -652 799 -632
rect 838 -652 848 -632
rect 852 -652 862 -632
rect 1709 -616 1719 -596
rect 1723 -616 1733 -596
rect 1768 -607 1778 -587
rect 1782 -607 1792 -587
rect 1824 -607 1834 -587
rect 1838 -607 1848 -587
rect 1879 -616 1889 -596
rect 1893 -616 1903 -596
rect 1938 -607 1948 -587
rect 1952 -607 1962 -587
rect 1994 -607 2004 -587
rect 2008 -607 2018 -587
rect 2049 -616 2059 -596
rect 2063 -616 2073 -596
rect 2108 -607 2118 -587
rect 2122 -607 2132 -587
rect 2164 -607 2174 -587
rect 2178 -607 2188 -587
rect 2219 -616 2229 -596
rect 2233 -616 2243 -596
rect 949 -688 959 -668
rect 963 -688 973 -668
rect 1005 -688 1015 -668
rect 1019 -688 1029 -668
rect 1103 -688 1113 -668
rect 1117 -688 1127 -668
rect 634 -734 644 -714
rect 648 -734 658 -714
rect 698 -737 708 -717
rect 712 -737 722 -717
rect 775 -734 785 -714
rect 789 -734 799 -714
rect 839 -737 849 -717
rect 853 -737 863 -717
rect 1103 -734 1113 -714
rect 1117 -734 1127 -714
rect 634 -833 644 -813
rect 648 -833 658 -813
rect 690 -833 700 -813
rect 704 -833 714 -813
rect 746 -833 756 -813
rect 760 -833 770 -813
rect 842 -832 852 -812
rect 856 -832 866 -812
rect 898 -832 908 -812
rect 912 -832 922 -812
rect 954 -832 964 -812
rect 968 -832 978 -812
rect 1010 -832 1020 -812
rect 1024 -832 1034 -812
rect 1134 -832 1144 -812
rect 1148 -832 1158 -812
rect 1190 -832 1200 -812
rect 1204 -832 1214 -812
rect 1246 -832 1256 -812
rect 1260 -832 1270 -812
rect 1302 -832 1312 -812
rect 1316 -832 1326 -812
rect 1416 -910 1426 -890
rect 1430 -910 1440 -890
rect 1472 -910 1482 -890
rect 1486 -910 1496 -890
rect 1527 -919 1537 -899
rect 1541 -919 1551 -899
<< psubstratepcontact >>
rect 462 461 466 465
rect 550 461 554 465
rect 573 461 577 465
rect 605 461 609 465
rect 637 461 641 465
rect 725 461 729 465
rect 748 461 752 465
rect 780 461 784 465
rect 812 461 816 465
rect 900 461 904 465
rect 923 461 927 465
rect 955 461 959 465
rect 987 461 991 465
rect 1075 461 1079 465
rect 1098 461 1102 465
rect 1130 461 1134 465
rect 1165 461 1169 465
rect 1253 461 1257 465
rect 1276 461 1280 465
rect 1308 461 1312 465
rect 1335 461 1339 465
rect 1423 461 1427 465
rect 1446 461 1450 465
rect 1478 461 1482 465
rect 1505 461 1509 465
rect 1593 461 1597 465
rect 1616 461 1620 465
rect 1648 461 1652 465
rect 1675 461 1679 465
rect 1763 461 1767 465
rect 1786 461 1790 465
rect 1818 461 1822 465
rect 462 310 466 314
rect 550 310 554 314
rect 573 310 577 314
rect 605 310 609 314
rect 637 310 641 314
rect 725 310 729 314
rect 748 310 752 314
rect 780 310 784 314
rect 812 310 816 314
rect 900 310 904 314
rect 923 310 927 314
rect 955 310 959 314
rect 987 310 991 314
rect 1075 310 1079 314
rect 1098 310 1102 314
rect 1130 310 1134 314
rect 2469 308 2473 312
rect 2501 308 2505 312
rect 2647 308 2651 312
rect 2679 308 2683 312
rect 2802 308 2806 312
rect 2834 308 2838 312
rect 2958 308 2962 312
rect 2990 308 2994 312
rect 2353 272 2357 276
rect 2385 272 2389 276
rect 1160 150 1164 154
rect 1248 150 1252 154
rect 1271 150 1275 154
rect 1303 150 1307 154
rect 1335 150 1339 154
rect 1423 150 1427 154
rect 1446 150 1450 154
rect 1478 150 1482 154
rect 1510 150 1514 154
rect 1598 150 1602 154
rect 1621 150 1625 154
rect 1653 150 1657 154
rect 1685 150 1689 154
rect 1773 150 1777 154
rect 1796 150 1800 154
rect 1828 150 1832 154
rect 558 137 562 141
rect 590 137 594 141
rect 616 137 620 141
rect 704 137 708 141
rect 727 137 731 141
rect 759 137 763 141
rect 786 137 790 141
rect 874 137 878 141
rect 897 137 901 141
rect 929 137 933 141
rect 2265 39 2269 43
rect 2353 39 2357 43
rect 2376 39 2380 43
rect 2408 39 2412 43
rect 2447 39 2451 43
rect 2535 39 2539 43
rect 2558 39 2562 43
rect 2590 39 2594 43
rect 2615 39 2619 43
rect 2708 39 2712 43
rect 2728 39 2732 43
rect 2760 39 2764 43
rect 2787 39 2791 43
rect 2875 39 2879 43
rect 2898 39 2902 43
rect 2930 39 2934 43
rect 2969 39 2973 43
rect 3057 39 3061 43
rect 3080 39 3084 43
rect 3112 39 3116 43
rect 3137 39 3141 43
rect 3230 39 3234 43
rect 3250 39 3254 43
rect 3282 39 3286 43
rect 558 -1 562 3
rect 590 -1 594 3
rect 616 -1 620 3
rect 704 -1 708 3
rect 727 -1 731 3
rect 759 -1 763 3
rect 786 -1 790 3
rect 874 -1 878 3
rect 897 -1 901 3
rect 929 -1 933 3
rect 982 -1 986 3
rect 1075 -1 1079 3
rect 1095 -1 1099 3
rect 1127 -1 1131 3
rect 1160 -1 1164 3
rect 1248 -1 1252 3
rect 1271 -1 1275 3
rect 1303 -1 1307 3
rect 1335 -1 1339 3
rect 1423 -1 1427 3
rect 1446 -1 1450 3
rect 1478 -1 1482 3
rect 1510 -1 1514 3
rect 1598 -1 1602 3
rect 1621 -1 1625 3
rect 1653 -1 1657 3
rect 1685 -1 1689 3
rect 1773 -1 1777 3
rect 1796 -1 1800 3
rect 1828 -1 1832 3
rect 2324 -43 2328 -39
rect 2356 -43 2360 -39
rect 2635 -40 2639 -36
rect 2667 -40 2671 -36
rect 2846 -43 2850 -39
rect 2878 -43 2882 -39
rect 3157 -40 3161 -36
rect 3189 -40 3193 -36
rect 2324 -125 2328 -121
rect 2356 -125 2360 -121
rect 2635 -122 2639 -118
rect 2667 -122 2671 -118
rect 2846 -125 2850 -121
rect 2878 -125 2882 -121
rect 3157 -122 3161 -118
rect 3189 -122 3193 -118
rect 505 -247 509 -243
rect 593 -247 597 -243
rect 616 -247 620 -243
rect 648 -247 652 -243
rect 680 -247 684 -243
rect 768 -247 772 -243
rect 791 -247 795 -243
rect 823 -247 827 -243
rect 855 -247 859 -243
rect 943 -247 947 -243
rect 966 -247 970 -243
rect 998 -247 1002 -243
rect 1030 -247 1034 -243
rect 1118 -247 1122 -243
rect 1141 -247 1145 -243
rect 1173 -247 1177 -243
rect 2265 -347 2269 -343
rect 2353 -347 2357 -343
rect 2376 -347 2380 -343
rect 2408 -347 2412 -343
rect 2447 -347 2451 -343
rect 2535 -347 2539 -343
rect 2558 -347 2562 -343
rect 2590 -347 2594 -343
rect 2615 -347 2619 -343
rect 2708 -347 2712 -343
rect 2728 -347 2732 -343
rect 2760 -347 2764 -343
rect 2787 -347 2791 -343
rect 2875 -347 2879 -343
rect 2898 -347 2902 -343
rect 2930 -347 2934 -343
rect 2969 -347 2973 -343
rect 3057 -347 3061 -343
rect 3080 -347 3084 -343
rect 3112 -347 3116 -343
rect 3137 -347 3141 -343
rect 3230 -347 3234 -343
rect 3250 -347 3254 -343
rect 3282 -347 3286 -343
rect 505 -398 509 -394
rect 593 -398 597 -394
rect 616 -398 620 -394
rect 648 -398 652 -394
rect 680 -398 684 -394
rect 768 -398 772 -394
rect 791 -398 795 -394
rect 823 -398 827 -394
rect 855 -398 859 -394
rect 943 -398 947 -394
rect 966 -398 970 -394
rect 998 -398 1002 -394
rect 1030 -398 1034 -394
rect 1118 -398 1122 -394
rect 1141 -398 1145 -394
rect 1173 -398 1177 -394
rect 2324 -429 2328 -425
rect 2356 -429 2360 -425
rect 2635 -426 2639 -422
rect 2667 -426 2671 -422
rect 2846 -429 2850 -425
rect 2878 -429 2882 -425
rect 3157 -426 3161 -422
rect 3189 -426 3193 -422
rect 628 -517 632 -513
rect 660 -517 664 -513
rect 769 -517 773 -513
rect 801 -517 805 -513
rect 2324 -511 2328 -507
rect 2356 -511 2360 -507
rect 2635 -508 2639 -504
rect 2667 -508 2671 -504
rect 2846 -511 2850 -507
rect 2878 -511 2882 -507
rect 3157 -508 3161 -504
rect 3189 -508 3193 -504
rect 628 -599 632 -595
rect 660 -599 664 -595
rect 769 -599 773 -595
rect 801 -599 805 -595
rect 913 -651 917 -647
rect 1113 -651 1117 -647
rect 1134 -651 1138 -647
rect 1166 -651 1170 -647
rect 628 -698 632 -694
rect 660 -698 664 -694
rect 769 -698 773 -694
rect 801 -698 805 -694
rect 1592 -709 1596 -705
rect 1680 -709 1684 -705
rect 1703 -709 1707 -705
rect 1735 -709 1739 -705
rect 1762 -709 1766 -705
rect 1850 -709 1854 -705
rect 1873 -709 1877 -705
rect 1905 -709 1909 -705
rect 1932 -709 1936 -705
rect 2020 -709 2024 -705
rect 2043 -709 2047 -705
rect 2075 -709 2079 -705
rect 2102 -709 2106 -705
rect 2190 -709 2194 -705
rect 2213 -709 2217 -705
rect 2245 -709 2249 -705
rect 628 -780 632 -776
rect 660 -780 664 -776
rect 1230 -755 1234 -751
rect 1485 -755 1489 -751
rect 769 -780 773 -776
rect 801 -780 805 -776
rect 943 -790 947 -786
rect 1031 -790 1035 -786
rect 1072 -794 1076 -790
rect 1165 -794 1169 -790
rect 628 -974 632 -970
rect 772 -974 776 -970
rect 836 -1012 840 -1008
rect 1036 -1012 1040 -1008
rect 1128 -1012 1132 -1008
rect 1328 -1012 1332 -1008
rect 1410 -1012 1414 -1008
rect 1498 -1012 1502 -1008
rect 1521 -1012 1525 -1008
rect 1553 -1012 1557 -1008
<< nsubstratencontact >>
rect 462 589 466 593
rect 550 589 554 593
rect 573 589 577 593
rect 605 589 609 593
rect 637 589 641 593
rect 725 589 729 593
rect 748 589 752 593
rect 780 589 784 593
rect 812 589 816 593
rect 900 589 904 593
rect 923 589 927 593
rect 955 589 959 593
rect 987 589 991 593
rect 1075 589 1079 593
rect 1098 589 1102 593
rect 1130 589 1134 593
rect 1165 589 1169 593
rect 1253 589 1257 593
rect 1276 589 1280 593
rect 1308 589 1312 593
rect 1335 589 1339 593
rect 1423 589 1427 593
rect 1446 589 1450 593
rect 1478 589 1482 593
rect 1505 589 1509 593
rect 1593 589 1597 593
rect 1616 589 1620 593
rect 1648 589 1652 593
rect 1675 589 1679 593
rect 1763 589 1767 593
rect 1786 589 1790 593
rect 1818 589 1822 593
rect 462 438 466 442
rect 550 438 554 442
rect 573 438 577 442
rect 605 438 609 442
rect 637 438 641 442
rect 725 438 729 442
rect 748 438 752 442
rect 780 438 784 442
rect 812 438 816 442
rect 900 438 904 442
rect 923 438 927 442
rect 955 438 959 442
rect 987 438 991 442
rect 1075 438 1079 442
rect 1098 438 1102 442
rect 1130 438 1134 442
rect 2469 380 2473 384
rect 2501 380 2505 384
rect 2647 380 2651 384
rect 2679 380 2683 384
rect 2802 380 2806 384
rect 2834 380 2838 384
rect 2958 380 2962 384
rect 2990 380 2994 384
rect 2353 344 2357 348
rect 2385 344 2389 348
rect 1160 278 1164 282
rect 1248 278 1252 282
rect 1271 278 1275 282
rect 1303 278 1307 282
rect 1335 278 1339 282
rect 1423 278 1427 282
rect 1446 278 1450 282
rect 1478 278 1482 282
rect 1510 278 1514 282
rect 1598 278 1602 282
rect 1621 278 1625 282
rect 1653 278 1657 282
rect 1685 278 1689 282
rect 1773 278 1777 282
rect 1796 278 1800 282
rect 1828 278 1832 282
rect 558 265 562 269
rect 590 265 594 269
rect 616 265 620 269
rect 704 265 708 269
rect 727 265 731 269
rect 759 265 763 269
rect 786 265 790 269
rect 874 265 878 269
rect 897 265 901 269
rect 929 265 933 269
rect 2265 171 2269 175
rect 2353 171 2357 175
rect 2376 171 2380 175
rect 2408 171 2412 175
rect 2447 171 2451 175
rect 2535 171 2539 175
rect 2558 171 2562 175
rect 2590 171 2594 175
rect 2640 171 2644 175
rect 2672 171 2676 175
rect 2728 171 2732 175
rect 2760 171 2764 175
rect 2787 171 2791 175
rect 2875 171 2879 175
rect 2898 171 2902 175
rect 2930 171 2934 175
rect 2969 171 2973 175
rect 3057 171 3061 175
rect 3080 171 3084 175
rect 3112 171 3116 175
rect 3162 171 3166 175
rect 3194 171 3198 175
rect 3250 171 3254 175
rect 3282 171 3286 175
rect 1007 131 1011 135
rect 1039 131 1043 135
rect 1095 131 1099 135
rect 1127 131 1131 135
rect 558 127 562 131
rect 590 127 594 131
rect 616 127 620 131
rect 704 127 708 131
rect 727 127 731 131
rect 759 127 763 131
rect 786 127 790 131
rect 874 127 878 131
rect 897 127 901 131
rect 929 127 933 131
rect 1160 127 1164 131
rect 1248 127 1252 131
rect 1271 127 1275 131
rect 1303 127 1307 131
rect 1335 127 1339 131
rect 1423 127 1427 131
rect 1446 127 1450 131
rect 1478 127 1482 131
rect 1510 127 1514 131
rect 1598 127 1602 131
rect 1621 127 1625 131
rect 1653 127 1657 131
rect 1685 127 1689 131
rect 1773 127 1777 131
rect 1796 127 1800 131
rect 1828 127 1832 131
rect 2324 29 2328 33
rect 2356 29 2360 33
rect 2635 32 2639 36
rect 2667 32 2671 36
rect 2846 29 2850 33
rect 2878 29 2882 33
rect 3157 32 3161 36
rect 3189 32 3193 36
rect 2324 -53 2328 -49
rect 2356 -53 2360 -49
rect 2635 -50 2639 -46
rect 2667 -50 2671 -46
rect 2846 -53 2850 -49
rect 2878 -53 2882 -49
rect 3157 -50 3161 -46
rect 3189 -50 3193 -46
rect 505 -119 509 -115
rect 593 -119 597 -115
rect 616 -119 620 -115
rect 648 -119 652 -115
rect 680 -119 684 -115
rect 768 -119 772 -115
rect 791 -119 795 -115
rect 823 -119 827 -115
rect 855 -119 859 -115
rect 943 -119 947 -115
rect 966 -119 970 -115
rect 998 -119 1002 -115
rect 1030 -119 1034 -115
rect 1118 -119 1122 -115
rect 1141 -119 1145 -115
rect 1173 -119 1177 -115
rect 2265 -215 2269 -211
rect 2353 -215 2357 -211
rect 2376 -215 2380 -211
rect 2408 -215 2412 -211
rect 2447 -215 2451 -211
rect 2535 -215 2539 -211
rect 2558 -215 2562 -211
rect 2590 -215 2594 -211
rect 2640 -215 2644 -211
rect 2672 -215 2676 -211
rect 2728 -215 2732 -211
rect 2760 -215 2764 -211
rect 2787 -215 2791 -211
rect 2875 -215 2879 -211
rect 2898 -215 2902 -211
rect 2930 -215 2934 -211
rect 2969 -215 2973 -211
rect 3057 -215 3061 -211
rect 3080 -215 3084 -211
rect 3112 -215 3116 -211
rect 3162 -215 3166 -211
rect 3194 -215 3198 -211
rect 3250 -215 3254 -211
rect 3282 -215 3286 -211
rect 505 -270 509 -266
rect 593 -270 597 -266
rect 616 -270 620 -266
rect 648 -270 652 -266
rect 680 -270 684 -266
rect 768 -270 772 -266
rect 791 -270 795 -266
rect 823 -270 827 -266
rect 855 -270 859 -266
rect 943 -270 947 -266
rect 966 -270 970 -266
rect 998 -270 1002 -266
rect 1030 -270 1034 -266
rect 1118 -270 1122 -266
rect 1141 -270 1145 -266
rect 1173 -270 1177 -266
rect 2324 -357 2328 -353
rect 2356 -357 2360 -353
rect 2635 -354 2639 -350
rect 2667 -354 2671 -350
rect 2846 -357 2850 -353
rect 2878 -357 2882 -353
rect 3157 -354 3161 -350
rect 3189 -354 3193 -350
rect 2324 -439 2328 -435
rect 2356 -439 2360 -435
rect 2635 -436 2639 -432
rect 2667 -436 2671 -432
rect 2846 -439 2850 -435
rect 2878 -439 2882 -435
rect 3157 -436 3161 -432
rect 3189 -436 3193 -432
rect 628 -445 632 -441
rect 660 -445 664 -441
rect 769 -445 773 -441
rect 801 -445 805 -441
rect 913 -445 917 -441
rect 1112 -445 1116 -441
rect 1134 -445 1138 -441
rect 1166 -445 1170 -441
rect 1230 -510 1234 -506
rect 1485 -510 1489 -506
rect 628 -527 632 -523
rect 660 -527 664 -523
rect 769 -527 773 -523
rect 801 -527 805 -523
rect 1592 -581 1596 -577
rect 1680 -581 1684 -577
rect 1703 -581 1707 -577
rect 1735 -581 1739 -577
rect 1762 -581 1766 -577
rect 1850 -581 1854 -577
rect 1873 -581 1877 -577
rect 1905 -581 1909 -577
rect 1932 -581 1936 -577
rect 2020 -581 2024 -577
rect 2043 -581 2047 -577
rect 2075 -581 2079 -577
rect 2102 -581 2106 -577
rect 2190 -581 2194 -577
rect 2213 -581 2217 -577
rect 2245 -581 2249 -577
rect 628 -626 632 -622
rect 660 -626 664 -622
rect 769 -626 773 -622
rect 801 -626 805 -622
rect 943 -662 947 -658
rect 1031 -662 1035 -658
rect 1097 -662 1101 -658
rect 1129 -662 1133 -658
rect 628 -708 632 -704
rect 660 -708 664 -704
rect 769 -708 773 -704
rect 801 -708 805 -704
rect 628 -807 632 -803
rect 772 -807 776 -803
rect 836 -806 840 -802
rect 1036 -806 1040 -802
rect 1128 -806 1132 -802
rect 1328 -806 1332 -802
rect 1410 -884 1414 -880
rect 1498 -884 1502 -880
rect 1521 -884 1525 -880
rect 1553 -884 1557 -880
<< polysilicon >>
rect 479 583 481 586
rect 535 583 537 586
rect 654 583 656 586
rect 710 583 712 586
rect 829 583 831 586
rect 885 583 887 586
rect 1004 583 1006 586
rect 1060 583 1062 586
rect 1182 583 1184 586
rect 1238 583 1240 586
rect 1352 583 1354 586
rect 1408 583 1410 586
rect 1522 583 1524 586
rect 1578 583 1580 586
rect 1692 583 1694 586
rect 1748 583 1750 586
rect 590 574 592 577
rect 479 554 481 563
rect 535 554 537 563
rect 765 574 767 577
rect 654 554 656 563
rect 710 554 712 563
rect 940 574 942 577
rect 829 554 831 563
rect 885 554 887 563
rect 1115 574 1117 577
rect 1004 554 1006 563
rect 1060 554 1062 563
rect 1293 574 1295 577
rect 1182 554 1184 563
rect 1238 554 1240 563
rect 1463 574 1465 577
rect 1352 554 1354 563
rect 1408 554 1410 563
rect 1633 574 1635 577
rect 1522 554 1524 563
rect 1578 554 1580 563
rect 1803 574 1805 577
rect 1692 554 1694 563
rect 1748 554 1750 563
rect 466 550 481 554
rect 522 550 537 554
rect 590 545 592 554
rect 641 550 656 554
rect 697 550 712 554
rect 765 545 767 554
rect 816 550 831 554
rect 872 550 887 554
rect 940 545 942 554
rect 991 550 1006 554
rect 1047 550 1062 554
rect 1115 545 1117 554
rect 1169 550 1184 554
rect 1225 550 1240 554
rect 1293 545 1295 554
rect 1339 550 1354 554
rect 1395 550 1410 554
rect 1463 545 1465 554
rect 1509 550 1524 554
rect 1565 550 1580 554
rect 1633 545 1635 554
rect 1679 550 1694 554
rect 1735 550 1750 554
rect 1803 545 1805 554
rect 575 543 592 545
rect 575 541 593 543
rect 750 543 767 545
rect 750 541 768 543
rect 925 543 942 545
rect 925 541 943 543
rect 1100 543 1117 545
rect 1100 541 1118 543
rect 1278 543 1295 545
rect 1278 541 1296 543
rect 1448 543 1465 545
rect 1448 541 1466 543
rect 1618 543 1635 545
rect 1618 541 1636 543
rect 1788 543 1805 545
rect 1788 541 1806 543
rect 589 538 593 541
rect 764 538 768 541
rect 939 538 943 541
rect 1114 538 1118 541
rect 1292 538 1296 541
rect 1462 538 1466 541
rect 1632 538 1636 541
rect 1802 538 1806 541
rect 494 534 509 538
rect 505 531 509 534
rect 669 534 684 538
rect 680 531 684 534
rect 589 515 593 518
rect 844 534 859 538
rect 855 531 859 534
rect 764 515 768 518
rect 1019 534 1034 538
rect 1030 531 1034 534
rect 939 515 943 518
rect 1197 534 1212 538
rect 1208 531 1212 534
rect 1114 515 1118 518
rect 1367 534 1382 538
rect 1378 531 1382 534
rect 1292 515 1296 518
rect 1537 534 1552 538
rect 1548 531 1552 534
rect 1462 515 1466 518
rect 1707 534 1722 538
rect 1718 531 1722 534
rect 1632 515 1636 518
rect 1802 515 1806 518
rect 505 508 509 511
rect 680 508 684 511
rect 855 508 859 511
rect 1030 508 1034 511
rect 1208 508 1212 511
rect 1378 508 1382 511
rect 1548 508 1552 511
rect 1718 508 1722 511
rect 494 494 509 498
rect 669 494 684 498
rect 844 494 859 498
rect 1019 494 1034 498
rect 1197 494 1212 498
rect 1367 494 1382 498
rect 1537 494 1552 498
rect 1707 494 1722 498
rect 505 491 509 494
rect 680 491 684 494
rect 855 491 859 494
rect 1030 491 1034 494
rect 1208 491 1212 494
rect 1378 491 1382 494
rect 1548 491 1552 494
rect 1718 491 1722 494
rect 505 468 509 471
rect 680 468 684 471
rect 855 468 859 471
rect 1030 468 1034 471
rect 1208 468 1212 471
rect 1378 468 1382 471
rect 1548 468 1552 471
rect 1718 468 1722 471
rect 479 432 481 435
rect 535 432 537 435
rect 654 432 656 435
rect 710 432 712 435
rect 829 432 831 435
rect 885 432 887 435
rect 1004 432 1006 435
rect 1060 432 1062 435
rect 590 423 592 426
rect 479 403 481 412
rect 535 403 537 412
rect 765 423 767 426
rect 654 403 656 412
rect 710 403 712 412
rect 940 423 942 426
rect 829 403 831 412
rect 885 403 887 412
rect 1115 423 1117 426
rect 1004 403 1006 412
rect 1060 403 1062 412
rect 466 399 481 403
rect 522 399 537 403
rect 590 394 592 403
rect 641 399 656 403
rect 697 399 712 403
rect 765 394 767 403
rect 816 399 831 403
rect 872 399 887 403
rect 940 394 942 403
rect 991 399 1006 403
rect 1047 399 1062 403
rect 1115 394 1117 403
rect 575 392 592 394
rect 575 390 593 392
rect 750 392 767 394
rect 750 390 768 392
rect 925 392 942 394
rect 925 390 943 392
rect 1100 392 1117 394
rect 1100 390 1118 392
rect 589 387 593 390
rect 764 387 768 390
rect 939 387 943 390
rect 1114 387 1118 390
rect 494 383 509 387
rect 505 380 509 383
rect 669 383 684 387
rect 680 380 684 383
rect 589 364 593 367
rect 844 383 859 387
rect 855 380 859 383
rect 764 364 768 367
rect 1019 383 1034 387
rect 1030 380 1034 383
rect 939 364 943 367
rect 2486 374 2488 377
rect 2549 374 2551 377
rect 2664 374 2666 377
rect 2727 374 2729 377
rect 2819 374 2821 377
rect 2882 374 2884 377
rect 2975 374 2977 377
rect 3038 374 3040 377
rect 1114 364 1118 367
rect 505 357 509 360
rect 680 357 684 360
rect 855 357 859 360
rect 1030 357 1034 360
rect 494 343 509 347
rect 669 343 684 347
rect 844 343 859 347
rect 1019 343 1034 347
rect 2486 345 2488 354
rect 2549 345 2551 354
rect 2664 345 2666 354
rect 2727 345 2729 354
rect 2819 345 2821 354
rect 2882 345 2884 354
rect 2975 345 2977 354
rect 3038 345 3040 354
rect 505 340 509 343
rect 680 340 684 343
rect 855 340 859 343
rect 1030 340 1034 343
rect 2471 343 2488 345
rect 2471 341 2489 343
rect 2534 341 2551 345
rect 2649 343 2666 345
rect 2649 341 2667 343
rect 2712 341 2729 345
rect 2804 343 2821 345
rect 2804 341 2822 343
rect 2867 341 2884 345
rect 2960 343 2977 345
rect 2960 341 2978 343
rect 3023 341 3040 345
rect 2370 338 2372 341
rect 2485 338 2489 341
rect 2663 338 2667 341
rect 2818 338 2822 341
rect 2974 338 2978 341
rect 505 317 509 320
rect 680 317 684 320
rect 855 317 859 320
rect 1030 317 1034 320
rect 2564 329 2568 332
rect 2370 309 2372 318
rect 2485 315 2489 318
rect 2355 307 2372 309
rect 2742 329 2746 332
rect 2663 315 2667 318
rect 2355 305 2373 307
rect 2564 306 2568 309
rect 2897 329 2901 332
rect 2818 315 2822 318
rect 2742 306 2746 309
rect 3053 329 3057 332
rect 2974 315 2978 318
rect 2897 306 2901 309
rect 3053 306 3057 309
rect 2369 302 2373 305
rect 2551 302 2568 306
rect 2729 302 2746 306
rect 2884 302 2901 306
rect 3040 302 3057 306
rect 2550 289 2552 292
rect 2728 289 2730 292
rect 2883 289 2885 292
rect 3039 289 3041 292
rect 2369 279 2373 282
rect 1177 272 1179 275
rect 1233 272 1235 275
rect 1352 272 1354 275
rect 1408 272 1410 275
rect 1527 272 1529 275
rect 1583 272 1585 275
rect 1702 272 1704 275
rect 1758 272 1760 275
rect 633 259 635 262
rect 689 259 691 262
rect 803 259 805 262
rect 859 259 861 262
rect 744 250 746 253
rect 633 230 635 239
rect 689 230 691 239
rect 914 250 916 253
rect 1288 263 1290 266
rect 803 230 805 239
rect 859 230 861 239
rect 1177 243 1179 252
rect 1233 243 1235 252
rect 1463 263 1465 266
rect 1352 243 1354 252
rect 1408 243 1410 252
rect 1638 263 1640 266
rect 1527 243 1529 252
rect 1583 243 1585 252
rect 1813 263 1815 266
rect 1702 243 1704 252
rect 1758 243 1760 252
rect 2550 260 2552 269
rect 2728 260 2730 269
rect 2883 260 2885 269
rect 3039 260 3041 269
rect 2535 256 2552 260
rect 2713 256 2730 260
rect 2868 256 2885 260
rect 3024 256 3041 260
rect 2565 244 2569 247
rect 2743 244 2747 247
rect 2898 244 2902 247
rect 3054 244 3058 247
rect 1164 239 1179 243
rect 1220 239 1235 243
rect 1288 234 1290 243
rect 1339 239 1354 243
rect 1395 239 1410 243
rect 1463 234 1465 243
rect 1514 239 1529 243
rect 1570 239 1585 243
rect 1638 234 1640 243
rect 1689 239 1704 243
rect 1745 239 1760 243
rect 1813 234 1815 243
rect 1273 232 1290 234
rect 1273 230 1291 232
rect 1448 232 1465 234
rect 1448 230 1466 232
rect 1623 232 1640 234
rect 1623 230 1641 232
rect 1798 232 1815 234
rect 1798 230 1816 232
rect 620 226 635 230
rect 676 226 691 230
rect 744 221 746 230
rect 790 226 805 230
rect 846 226 861 230
rect 914 221 916 230
rect 1287 227 1291 230
rect 1462 227 1466 230
rect 1637 227 1641 230
rect 1812 227 1816 230
rect 1192 223 1207 227
rect 729 219 746 221
rect 729 217 747 219
rect 899 219 916 221
rect 1203 220 1207 223
rect 899 217 917 219
rect 743 214 747 217
rect 913 214 917 217
rect 648 210 663 214
rect 659 207 663 210
rect 575 203 577 206
rect 818 210 833 214
rect 829 207 833 210
rect 743 191 747 194
rect 1367 223 1382 227
rect 1378 220 1382 223
rect 1287 204 1291 207
rect 1542 223 1557 227
rect 1553 220 1557 223
rect 1462 204 1466 207
rect 1717 223 1732 227
rect 1728 220 1732 223
rect 1637 204 1641 207
rect 2565 221 2569 224
rect 2743 221 2747 224
rect 2898 221 2902 224
rect 3054 221 3058 224
rect 2552 217 2569 221
rect 2730 217 2747 221
rect 2885 217 2902 221
rect 3041 217 3058 221
rect 1812 204 1816 207
rect 1203 197 1207 200
rect 1378 197 1382 200
rect 1553 197 1557 200
rect 1728 197 1732 200
rect 913 191 917 194
rect 659 184 663 187
rect 829 184 833 187
rect 1192 183 1207 187
rect 1367 183 1382 187
rect 1542 183 1557 187
rect 1717 183 1732 187
rect 575 174 577 183
rect 1203 180 1207 183
rect 1378 180 1382 183
rect 1553 180 1557 183
rect 1728 180 1732 183
rect 560 172 577 174
rect 560 170 578 172
rect 648 170 663 174
rect 818 170 833 174
rect 574 167 578 170
rect 659 167 663 170
rect 829 167 833 170
rect 2657 165 2659 168
rect 3179 165 3181 168
rect 2282 161 2284 164
rect 2338 161 2340 164
rect 2464 161 2466 164
rect 2520 161 2522 164
rect 1203 157 1207 160
rect 1378 157 1382 160
rect 1553 157 1557 160
rect 1728 157 1732 160
rect 574 144 578 147
rect 659 144 663 147
rect 829 144 833 147
rect 2393 152 2395 155
rect 2282 132 2284 141
rect 2338 132 2340 141
rect 2575 152 2577 155
rect 2464 132 2466 141
rect 2520 132 2522 141
rect 2804 161 2806 164
rect 2860 161 2862 164
rect 2986 161 2988 164
rect 3042 161 3044 164
rect 2657 136 2659 145
rect 2915 152 2917 155
rect 2644 132 2659 136
rect 2804 132 2806 141
rect 2860 132 2862 141
rect 3097 152 3099 155
rect 2986 132 2988 141
rect 3042 132 3044 141
rect 3179 136 3181 145
rect 3166 132 3181 136
rect 1024 125 1026 128
rect 2269 128 2284 132
rect 2325 128 2340 132
rect 633 121 635 124
rect 689 121 691 124
rect 803 121 805 124
rect 859 121 861 124
rect 744 112 746 115
rect 633 92 635 101
rect 689 92 691 101
rect 914 112 916 115
rect 803 92 805 101
rect 859 92 861 101
rect 1177 121 1179 124
rect 1233 121 1235 124
rect 1352 121 1354 124
rect 1408 121 1410 124
rect 1527 121 1529 124
rect 1583 121 1585 124
rect 1702 121 1704 124
rect 1758 121 1760 124
rect 2393 123 2395 132
rect 2451 128 2466 132
rect 2507 128 2522 132
rect 2575 123 2577 132
rect 2791 128 2806 132
rect 2847 128 2862 132
rect 2915 123 2917 132
rect 2973 128 2988 132
rect 3029 128 3044 132
rect 3097 123 3099 132
rect 1024 96 1026 105
rect 1288 112 1290 115
rect 1011 92 1026 96
rect 1177 92 1179 101
rect 1233 92 1235 101
rect 1463 112 1465 115
rect 1352 92 1354 101
rect 1408 92 1410 101
rect 1638 112 1640 115
rect 1527 92 1529 101
rect 1583 92 1585 101
rect 2378 121 2395 123
rect 2378 119 2396 121
rect 2560 121 2577 123
rect 2560 119 2578 121
rect 2657 119 2659 122
rect 2900 121 2917 123
rect 2900 119 2918 121
rect 3082 121 3099 123
rect 3082 119 3100 121
rect 3179 119 3181 122
rect 2392 116 2396 119
rect 2574 116 2578 119
rect 1813 112 1815 115
rect 2297 112 2312 116
rect 1702 92 1704 101
rect 1758 92 1760 101
rect 2308 109 2312 112
rect 620 88 635 92
rect 676 88 691 92
rect 744 83 746 92
rect 790 88 805 92
rect 846 88 861 92
rect 914 83 916 92
rect 1164 88 1179 92
rect 1220 88 1235 92
rect 1288 83 1290 92
rect 1339 88 1354 92
rect 1395 88 1410 92
rect 1463 83 1465 92
rect 1514 88 1529 92
rect 1570 88 1585 92
rect 1638 83 1640 92
rect 1689 88 1704 92
rect 1745 88 1760 92
rect 1813 83 1815 92
rect 2479 112 2494 116
rect 2490 109 2494 112
rect 2392 93 2396 96
rect 2914 116 2918 119
rect 3096 116 3100 119
rect 2745 112 2747 115
rect 2819 112 2834 116
rect 2574 93 2578 96
rect 2657 90 2659 99
rect 2830 109 2834 112
rect 2308 86 2312 89
rect 2490 86 2494 89
rect 2644 86 2659 90
rect 2745 83 2747 92
rect 3001 112 3016 116
rect 3012 109 3016 112
rect 2914 93 2918 96
rect 3267 112 3269 115
rect 3096 93 3100 96
rect 3179 90 3181 99
rect 2830 86 2834 89
rect 3012 86 3016 89
rect 3166 86 3181 90
rect 3267 83 3269 92
rect 729 81 746 83
rect 729 79 747 81
rect 899 81 916 83
rect 899 79 917 81
rect 1024 79 1026 82
rect 1273 81 1290 83
rect 1273 79 1291 81
rect 1448 81 1465 83
rect 1448 79 1466 81
rect 1623 81 1640 83
rect 1623 79 1641 81
rect 1798 81 1815 83
rect 1798 79 1816 81
rect 2730 81 2747 83
rect 2730 79 2748 81
rect 3252 81 3269 83
rect 3252 79 3270 81
rect 743 76 747 79
rect 913 76 917 79
rect 648 72 663 76
rect 659 69 663 72
rect 575 65 577 68
rect 818 72 833 76
rect 829 69 833 72
rect 743 53 747 56
rect 1287 76 1291 79
rect 1462 76 1466 79
rect 1637 76 1641 79
rect 1812 76 1816 79
rect 2744 76 2748 79
rect 3266 76 3270 79
rect 1112 72 1114 75
rect 1192 72 1207 76
rect 913 53 917 56
rect 1024 50 1026 59
rect 1203 69 1207 72
rect 659 46 663 49
rect 829 46 833 49
rect 1011 46 1026 50
rect 575 36 577 45
rect 1112 43 1114 52
rect 1367 72 1382 76
rect 1378 69 1382 72
rect 1287 53 1291 56
rect 1542 72 1557 76
rect 1553 69 1557 72
rect 1462 53 1466 56
rect 1717 72 1732 76
rect 1728 69 1732 72
rect 1637 53 1641 56
rect 2297 72 2312 76
rect 2479 72 2494 76
rect 2646 73 2650 76
rect 2697 73 2701 76
rect 2308 69 2312 72
rect 2490 69 2494 72
rect 1812 53 1816 56
rect 2819 72 2834 76
rect 3001 72 3016 76
rect 3168 73 3172 76
rect 3219 73 3223 76
rect 2830 69 2834 72
rect 3012 69 3016 72
rect 2744 53 2748 56
rect 2646 50 2650 53
rect 2697 50 2701 53
rect 1203 46 1207 49
rect 1378 46 1382 49
rect 1553 46 1557 49
rect 1728 46 1732 49
rect 2308 46 2312 49
rect 2490 46 2494 49
rect 2633 46 2650 50
rect 2684 46 2701 50
rect 3266 53 3270 56
rect 3168 50 3172 53
rect 3219 50 3223 53
rect 2830 46 2834 49
rect 3012 46 3016 49
rect 3155 46 3172 50
rect 3206 46 3223 50
rect 1097 41 1114 43
rect 1097 39 1115 41
rect 1111 36 1115 39
rect 560 34 577 36
rect 560 32 578 34
rect 648 32 663 36
rect 818 32 833 36
rect 1013 33 1017 36
rect 1064 33 1068 36
rect 574 29 578 32
rect 659 29 663 32
rect 829 29 833 32
rect 1192 32 1207 36
rect 1367 32 1382 36
rect 1542 32 1557 36
rect 1717 32 1732 36
rect 1203 29 1207 32
rect 1378 29 1382 32
rect 1553 29 1557 32
rect 1728 29 1732 32
rect 1111 13 1115 16
rect 1013 10 1017 13
rect 1064 10 1068 13
rect 574 6 578 9
rect 659 6 663 9
rect 829 6 833 9
rect 1000 6 1017 10
rect 1051 6 1068 10
rect 2652 26 2654 29
rect 2715 26 2717 29
rect 3174 26 3176 29
rect 3237 26 3239 29
rect 2341 23 2343 26
rect 2404 23 2406 26
rect 1203 6 1207 9
rect 1378 6 1382 9
rect 1553 6 1557 9
rect 1728 6 1732 9
rect 2863 23 2865 26
rect 2926 23 2928 26
rect 2341 -6 2343 3
rect 2404 -6 2406 3
rect 2652 -3 2654 6
rect 2715 -3 2717 6
rect 2326 -8 2343 -6
rect 2326 -10 2344 -8
rect 2389 -10 2406 -6
rect 2637 -5 2654 -3
rect 2637 -7 2655 -5
rect 2700 -7 2717 -3
rect 2863 -6 2865 3
rect 2926 -6 2928 3
rect 3174 -3 3176 6
rect 3237 -3 3239 6
rect 2651 -10 2655 -7
rect 2848 -8 2865 -6
rect 2848 -10 2866 -8
rect 2911 -10 2928 -6
rect 3159 -5 3176 -3
rect 3159 -7 3177 -5
rect 3222 -7 3239 -3
rect 3173 -10 3177 -7
rect 2340 -13 2344 -10
rect 2419 -22 2423 -19
rect 2340 -36 2344 -33
rect 2862 -13 2866 -10
rect 2730 -19 2734 -16
rect 2651 -33 2655 -30
rect 2941 -22 2945 -19
rect 2862 -36 2866 -33
rect 2730 -42 2734 -39
rect 2419 -45 2423 -42
rect 2406 -49 2423 -45
rect 2717 -46 2734 -42
rect 3252 -19 3256 -16
rect 3173 -33 3177 -30
rect 3252 -42 3256 -39
rect 2941 -45 2945 -42
rect 2928 -49 2945 -45
rect 3239 -46 3256 -42
rect 2652 -56 2654 -53
rect 3174 -56 3176 -53
rect 2341 -59 2343 -56
rect 2405 -62 2407 -59
rect 2341 -88 2343 -79
rect 2716 -59 2718 -56
rect 2863 -59 2865 -56
rect 2326 -90 2343 -88
rect 2326 -92 2344 -90
rect 2405 -91 2407 -82
rect 2652 -85 2654 -76
rect 2927 -62 2929 -59
rect 2637 -87 2654 -85
rect 2637 -89 2655 -87
rect 2716 -88 2718 -79
rect 2863 -88 2865 -79
rect 3238 -59 3240 -56
rect 2340 -95 2344 -92
rect 2390 -95 2407 -91
rect 2651 -92 2655 -89
rect 2701 -92 2718 -88
rect 2848 -90 2865 -88
rect 2848 -92 2866 -90
rect 2927 -91 2929 -82
rect 3174 -85 3176 -76
rect 3159 -87 3176 -85
rect 3159 -89 3177 -87
rect 3238 -88 3240 -79
rect 2420 -107 2424 -104
rect 2340 -118 2344 -115
rect 522 -125 524 -122
rect 578 -125 580 -122
rect 697 -125 699 -122
rect 753 -125 755 -122
rect 872 -125 874 -122
rect 928 -125 930 -122
rect 1047 -125 1049 -122
rect 1103 -125 1105 -122
rect 633 -134 635 -131
rect 522 -154 524 -145
rect 578 -154 580 -145
rect 808 -134 810 -131
rect 697 -154 699 -145
rect 753 -154 755 -145
rect 983 -134 985 -131
rect 872 -154 874 -145
rect 928 -154 930 -145
rect 2862 -95 2866 -92
rect 2912 -95 2929 -91
rect 3173 -92 3177 -89
rect 3223 -92 3240 -88
rect 2731 -104 2735 -101
rect 2651 -115 2655 -112
rect 2942 -107 2946 -104
rect 2862 -118 2866 -115
rect 2731 -127 2735 -124
rect 3253 -104 3257 -101
rect 3173 -115 3177 -112
rect 3253 -127 3257 -124
rect 2420 -130 2424 -127
rect 1158 -134 1160 -131
rect 2407 -134 2424 -130
rect 2718 -131 2735 -127
rect 2942 -130 2946 -127
rect 2929 -134 2946 -130
rect 3240 -131 3257 -127
rect 1047 -154 1049 -145
rect 1103 -154 1105 -145
rect 509 -158 524 -154
rect 565 -158 580 -154
rect 633 -163 635 -154
rect 684 -158 699 -154
rect 740 -158 755 -154
rect 808 -163 810 -154
rect 859 -158 874 -154
rect 915 -158 930 -154
rect 983 -163 985 -154
rect 1034 -158 1049 -154
rect 1090 -158 1105 -154
rect 1158 -163 1160 -154
rect 618 -165 635 -163
rect 618 -167 636 -165
rect 793 -165 810 -163
rect 793 -167 811 -165
rect 968 -165 985 -163
rect 968 -167 986 -165
rect 1143 -165 1160 -163
rect 1143 -167 1161 -165
rect 632 -170 636 -167
rect 807 -170 811 -167
rect 982 -170 986 -167
rect 1157 -170 1161 -167
rect 537 -174 552 -170
rect 548 -177 552 -174
rect 712 -174 727 -170
rect 723 -177 727 -174
rect 632 -193 636 -190
rect 887 -174 902 -170
rect 898 -177 902 -174
rect 807 -193 811 -190
rect 1062 -174 1077 -170
rect 1073 -177 1077 -174
rect 982 -193 986 -190
rect 1157 -193 1161 -190
rect 548 -200 552 -197
rect 723 -200 727 -197
rect 898 -200 902 -197
rect 1073 -200 1077 -197
rect 537 -214 552 -210
rect 712 -214 727 -210
rect 887 -214 902 -210
rect 1062 -214 1077 -210
rect 548 -217 552 -214
rect 723 -217 727 -214
rect 898 -217 902 -214
rect 1073 -217 1077 -214
rect 2657 -221 2659 -218
rect 3179 -221 3181 -218
rect 2282 -225 2284 -222
rect 2338 -225 2340 -222
rect 2464 -225 2466 -222
rect 2520 -225 2522 -222
rect 548 -240 552 -237
rect 723 -240 727 -237
rect 898 -240 902 -237
rect 1073 -240 1077 -237
rect 2393 -234 2395 -231
rect 2282 -254 2284 -245
rect 2338 -254 2340 -245
rect 2575 -234 2577 -231
rect 2464 -254 2466 -245
rect 2520 -254 2522 -245
rect 2804 -225 2806 -222
rect 2860 -225 2862 -222
rect 2986 -225 2988 -222
rect 3042 -225 3044 -222
rect 2657 -250 2659 -241
rect 2915 -234 2917 -231
rect 2644 -254 2659 -250
rect 2804 -254 2806 -245
rect 2860 -254 2862 -245
rect 3097 -234 3099 -231
rect 2986 -254 2988 -245
rect 3042 -254 3044 -245
rect 3179 -250 3181 -241
rect 3166 -254 3181 -250
rect 2269 -258 2284 -254
rect 2325 -258 2340 -254
rect 2393 -263 2395 -254
rect 2451 -258 2466 -254
rect 2507 -258 2522 -254
rect 2575 -263 2577 -254
rect 2791 -258 2806 -254
rect 2847 -258 2862 -254
rect 2915 -263 2917 -254
rect 2973 -258 2988 -254
rect 3029 -258 3044 -254
rect 3097 -263 3099 -254
rect 2378 -265 2395 -263
rect 2378 -267 2396 -265
rect 2560 -265 2577 -263
rect 2560 -267 2578 -265
rect 2657 -267 2659 -264
rect 2900 -265 2917 -263
rect 2900 -267 2918 -265
rect 3082 -265 3099 -263
rect 3082 -267 3100 -265
rect 3179 -267 3181 -264
rect 2392 -270 2396 -267
rect 2574 -270 2578 -267
rect 522 -276 524 -273
rect 578 -276 580 -273
rect 697 -276 699 -273
rect 753 -276 755 -273
rect 872 -276 874 -273
rect 928 -276 930 -273
rect 1047 -276 1049 -273
rect 1103 -276 1105 -273
rect 2297 -274 2312 -270
rect 633 -285 635 -282
rect 522 -305 524 -296
rect 578 -305 580 -296
rect 808 -285 810 -282
rect 697 -305 699 -296
rect 753 -305 755 -296
rect 983 -285 985 -282
rect 872 -305 874 -296
rect 928 -305 930 -296
rect 2308 -277 2312 -274
rect 1158 -285 1160 -282
rect 1047 -305 1049 -296
rect 1103 -305 1105 -296
rect 2479 -274 2494 -270
rect 2490 -277 2494 -274
rect 2392 -293 2396 -290
rect 2914 -270 2918 -267
rect 3096 -270 3100 -267
rect 2745 -274 2747 -271
rect 2819 -274 2834 -270
rect 2574 -293 2578 -290
rect 2657 -296 2659 -287
rect 2830 -277 2834 -274
rect 2308 -300 2312 -297
rect 2490 -300 2494 -297
rect 2644 -300 2659 -296
rect 2745 -303 2747 -294
rect 3001 -274 3016 -270
rect 3012 -277 3016 -274
rect 2914 -293 2918 -290
rect 3267 -274 3269 -271
rect 3096 -293 3100 -290
rect 3179 -296 3181 -287
rect 2830 -300 2834 -297
rect 3012 -300 3016 -297
rect 3166 -300 3181 -296
rect 3267 -303 3269 -294
rect 509 -309 524 -305
rect 565 -309 580 -305
rect 633 -314 635 -305
rect 684 -309 699 -305
rect 740 -309 755 -305
rect 808 -314 810 -305
rect 859 -309 874 -305
rect 915 -309 930 -305
rect 983 -314 985 -305
rect 1034 -309 1049 -305
rect 1090 -309 1105 -305
rect 1158 -314 1160 -305
rect 2730 -305 2747 -303
rect 2730 -307 2748 -305
rect 3252 -305 3269 -303
rect 3252 -307 3270 -305
rect 2744 -310 2748 -307
rect 3266 -310 3270 -307
rect 2297 -314 2312 -310
rect 2479 -314 2494 -310
rect 2646 -313 2650 -310
rect 2697 -313 2701 -310
rect 618 -316 635 -314
rect 618 -318 636 -316
rect 793 -316 810 -314
rect 793 -318 811 -316
rect 968 -316 985 -314
rect 968 -318 986 -316
rect 1143 -316 1160 -314
rect 1143 -318 1161 -316
rect 2308 -317 2312 -314
rect 2490 -317 2494 -314
rect 632 -321 636 -318
rect 807 -321 811 -318
rect 982 -321 986 -318
rect 1157 -321 1161 -318
rect 537 -325 552 -321
rect 548 -328 552 -325
rect 712 -325 727 -321
rect 723 -328 727 -325
rect 632 -344 636 -341
rect 887 -325 902 -321
rect 898 -328 902 -325
rect 807 -344 811 -341
rect 1062 -325 1077 -321
rect 1073 -328 1077 -325
rect 982 -344 986 -341
rect 2819 -314 2834 -310
rect 3001 -314 3016 -310
rect 3168 -313 3172 -310
rect 3219 -313 3223 -310
rect 2830 -317 2834 -314
rect 3012 -317 3016 -314
rect 2744 -333 2748 -330
rect 2646 -336 2650 -333
rect 2697 -336 2701 -333
rect 2308 -340 2312 -337
rect 2490 -340 2494 -337
rect 2633 -340 2650 -336
rect 2684 -340 2701 -336
rect 3266 -333 3270 -330
rect 3168 -336 3172 -333
rect 3219 -336 3223 -333
rect 2830 -340 2834 -337
rect 3012 -340 3016 -337
rect 3155 -340 3172 -336
rect 3206 -340 3223 -336
rect 1157 -344 1161 -341
rect 548 -351 552 -348
rect 723 -351 727 -348
rect 898 -351 902 -348
rect 1073 -351 1077 -348
rect 2652 -360 2654 -357
rect 2715 -360 2717 -357
rect 3174 -360 3176 -357
rect 3237 -360 3239 -357
rect 537 -365 552 -361
rect 712 -365 727 -361
rect 887 -365 902 -361
rect 1062 -365 1077 -361
rect 2341 -363 2343 -360
rect 2404 -363 2406 -360
rect 548 -368 552 -365
rect 723 -368 727 -365
rect 898 -368 902 -365
rect 1073 -368 1077 -365
rect 2863 -363 2865 -360
rect 2926 -363 2928 -360
rect 548 -391 552 -388
rect 723 -391 727 -388
rect 898 -391 902 -388
rect 1073 -391 1077 -388
rect 2341 -392 2343 -383
rect 2404 -392 2406 -383
rect 2652 -389 2654 -380
rect 2715 -389 2717 -380
rect 2326 -394 2343 -392
rect 2326 -396 2344 -394
rect 2389 -396 2406 -392
rect 2637 -391 2654 -389
rect 2637 -393 2655 -391
rect 2700 -393 2717 -389
rect 2863 -392 2865 -383
rect 2926 -392 2928 -383
rect 3174 -389 3176 -380
rect 3237 -389 3239 -380
rect 2651 -396 2655 -393
rect 2848 -394 2865 -392
rect 2848 -396 2866 -394
rect 2911 -396 2928 -392
rect 3159 -391 3176 -389
rect 3159 -393 3177 -391
rect 3222 -393 3239 -389
rect 3173 -396 3177 -393
rect 2340 -399 2344 -396
rect 2419 -408 2423 -405
rect 2340 -422 2344 -419
rect 2862 -399 2866 -396
rect 2730 -405 2734 -402
rect 2651 -419 2655 -416
rect 2941 -408 2945 -405
rect 2862 -422 2866 -419
rect 2730 -428 2734 -425
rect 2419 -431 2423 -428
rect 2406 -435 2423 -431
rect 2717 -432 2734 -428
rect 3252 -405 3256 -402
rect 3173 -419 3177 -416
rect 3252 -428 3256 -425
rect 2941 -431 2945 -428
rect 2928 -435 2945 -431
rect 3239 -432 3256 -428
rect 2652 -442 2654 -439
rect 3174 -442 3176 -439
rect 2341 -445 2343 -442
rect 645 -451 647 -448
rect 708 -451 710 -448
rect 786 -451 788 -448
rect 849 -451 851 -448
rect 930 -451 932 -448
rect 986 -451 988 -448
rect 1042 -451 1044 -448
rect 1098 -451 1100 -448
rect 1150 -460 1152 -457
rect 645 -480 647 -471
rect 708 -480 710 -471
rect 786 -480 788 -471
rect 849 -480 851 -471
rect 930 -480 932 -471
rect 986 -480 988 -471
rect 1042 -480 1044 -471
rect 1098 -480 1100 -471
rect 2405 -448 2407 -445
rect 2341 -474 2343 -465
rect 2716 -445 2718 -442
rect 2863 -445 2865 -442
rect 2326 -476 2343 -474
rect 2326 -478 2344 -476
rect 2405 -477 2407 -468
rect 2652 -471 2654 -462
rect 2927 -448 2929 -445
rect 2637 -473 2654 -471
rect 2637 -475 2655 -473
rect 2716 -474 2718 -465
rect 2863 -474 2865 -465
rect 3238 -445 3240 -442
rect 630 -482 647 -480
rect 630 -484 648 -482
rect 693 -484 710 -480
rect 771 -482 788 -480
rect 771 -484 789 -482
rect 834 -484 851 -480
rect 917 -484 932 -480
rect 973 -484 988 -480
rect 1029 -484 1044 -480
rect 1085 -484 1100 -480
rect 644 -487 648 -484
rect 785 -487 789 -484
rect 723 -496 727 -493
rect 644 -510 648 -507
rect 1150 -489 1152 -480
rect 2340 -481 2344 -478
rect 2390 -481 2407 -477
rect 2651 -478 2655 -475
rect 2701 -478 2718 -474
rect 2848 -476 2865 -474
rect 2848 -478 2866 -476
rect 2927 -477 2929 -468
rect 3174 -471 3176 -462
rect 3159 -473 3176 -471
rect 3159 -475 3177 -473
rect 3238 -474 3240 -465
rect 1135 -491 1152 -489
rect 1135 -493 1153 -491
rect 864 -496 868 -493
rect 1149 -496 1153 -493
rect 785 -510 789 -507
rect 723 -519 727 -516
rect 945 -500 960 -496
rect 956 -503 960 -500
rect 864 -519 868 -516
rect 710 -523 727 -519
rect 851 -523 868 -519
rect 2420 -493 2424 -490
rect 2340 -504 2344 -501
rect 2862 -481 2866 -478
rect 2912 -481 2929 -477
rect 3173 -478 3177 -475
rect 3223 -478 3240 -474
rect 2731 -490 2735 -487
rect 2651 -501 2655 -498
rect 2942 -493 2946 -490
rect 2862 -504 2866 -501
rect 2731 -513 2735 -510
rect 3253 -490 3257 -487
rect 3173 -501 3177 -498
rect 3253 -513 3257 -510
rect 1247 -516 1249 -513
rect 1303 -516 1305 -513
rect 1359 -516 1361 -513
rect 1415 -516 1417 -513
rect 1470 -516 1472 -513
rect 2420 -516 2424 -513
rect 1149 -519 1153 -516
rect 956 -526 960 -523
rect 645 -533 647 -530
rect 786 -533 788 -530
rect 709 -536 711 -533
rect 645 -562 647 -553
rect 850 -536 852 -533
rect 2407 -520 2424 -516
rect 2718 -517 2735 -513
rect 2942 -516 2946 -513
rect 2929 -520 2946 -516
rect 3240 -517 3257 -513
rect 630 -564 647 -562
rect 630 -566 648 -564
rect 709 -565 711 -556
rect 786 -562 788 -553
rect 945 -540 960 -536
rect 956 -543 960 -540
rect 644 -569 648 -566
rect 694 -569 711 -565
rect 771 -564 788 -562
rect 771 -566 789 -564
rect 850 -565 852 -556
rect 1247 -545 1249 -536
rect 1303 -545 1305 -536
rect 1359 -545 1361 -536
rect 1415 -545 1417 -536
rect 1470 -545 1472 -536
rect 1234 -549 1249 -545
rect 1290 -549 1305 -545
rect 1346 -549 1361 -545
rect 1402 -549 1417 -545
rect 1457 -549 1472 -545
rect 785 -569 789 -566
rect 835 -569 852 -565
rect 956 -566 960 -563
rect 1262 -565 1277 -561
rect 1273 -568 1277 -565
rect 724 -581 728 -578
rect 644 -592 648 -589
rect 865 -581 869 -578
rect 945 -580 960 -576
rect 785 -592 789 -589
rect 956 -583 960 -580
rect 724 -604 728 -601
rect 865 -604 869 -601
rect 1609 -587 1611 -584
rect 1665 -587 1667 -584
rect 1779 -587 1781 -584
rect 1835 -587 1837 -584
rect 1949 -587 1951 -584
rect 2005 -587 2007 -584
rect 2119 -587 2121 -584
rect 2175 -587 2177 -584
rect 1273 -591 1277 -588
rect 711 -608 728 -604
rect 852 -608 869 -604
rect 956 -606 960 -603
rect 1262 -605 1277 -601
rect 1273 -608 1277 -605
rect 1720 -596 1722 -593
rect 945 -619 960 -615
rect 956 -622 960 -619
rect 645 -632 647 -629
rect 708 -632 710 -629
rect 786 -632 788 -629
rect 849 -632 851 -629
rect 1609 -616 1611 -607
rect 1665 -616 1667 -607
rect 1890 -596 1892 -593
rect 1779 -616 1781 -607
rect 1835 -616 1837 -607
rect 2060 -596 2062 -593
rect 1949 -616 1951 -607
rect 2005 -616 2007 -607
rect 2230 -596 2232 -593
rect 2119 -616 2121 -607
rect 2175 -616 2177 -607
rect 1596 -620 1611 -616
rect 1652 -620 1667 -616
rect 1720 -625 1722 -616
rect 1766 -620 1781 -616
rect 1822 -620 1837 -616
rect 1890 -625 1892 -616
rect 1936 -620 1951 -616
rect 1992 -620 2007 -616
rect 2060 -625 2062 -616
rect 2106 -620 2121 -616
rect 2162 -620 2177 -616
rect 2230 -625 2232 -616
rect 1273 -631 1277 -628
rect 1705 -627 1722 -625
rect 1705 -629 1723 -627
rect 1875 -627 1892 -625
rect 1875 -629 1893 -627
rect 2045 -627 2062 -625
rect 2045 -629 2063 -627
rect 2215 -627 2232 -625
rect 2215 -629 2233 -627
rect 1719 -632 1723 -629
rect 1889 -632 1893 -629
rect 2059 -632 2063 -629
rect 2229 -632 2233 -629
rect 1624 -636 1639 -632
rect 1635 -639 1639 -636
rect 956 -645 960 -642
rect 1262 -645 1277 -641
rect 1273 -648 1277 -645
rect 645 -661 647 -652
rect 708 -661 710 -652
rect 786 -661 788 -652
rect 849 -661 851 -652
rect 630 -663 647 -661
rect 630 -665 648 -663
rect 693 -665 710 -661
rect 771 -663 788 -661
rect 771 -665 789 -663
rect 834 -665 851 -661
rect 644 -668 648 -665
rect 785 -668 789 -665
rect 960 -668 962 -665
rect 1016 -668 1018 -665
rect 1114 -668 1116 -665
rect 1794 -636 1809 -632
rect 1805 -639 1809 -636
rect 1719 -655 1723 -652
rect 1964 -636 1979 -632
rect 1975 -639 1979 -636
rect 1889 -655 1893 -652
rect 2134 -636 2149 -632
rect 2145 -639 2149 -636
rect 2059 -655 2063 -652
rect 2229 -655 2233 -652
rect 1635 -662 1639 -659
rect 1805 -662 1809 -659
rect 1975 -662 1979 -659
rect 2145 -662 2149 -659
rect 723 -677 727 -674
rect 644 -691 648 -688
rect 864 -677 868 -674
rect 785 -691 789 -688
rect 723 -700 727 -697
rect 1273 -671 1277 -668
rect 1624 -676 1639 -672
rect 1794 -676 1809 -672
rect 1964 -676 1979 -672
rect 2134 -676 2149 -672
rect 1635 -679 1639 -676
rect 1805 -679 1809 -676
rect 1975 -679 1979 -676
rect 2145 -679 2149 -676
rect 1262 -684 1277 -680
rect 1273 -687 1277 -684
rect 960 -697 962 -688
rect 1016 -697 1018 -688
rect 1114 -697 1116 -688
rect 864 -700 868 -697
rect 710 -704 727 -700
rect 851 -704 868 -700
rect 947 -701 962 -697
rect 1003 -701 1018 -697
rect 1101 -701 1116 -697
rect 1635 -702 1639 -699
rect 1805 -702 1809 -699
rect 1975 -702 1979 -699
rect 2145 -702 2149 -699
rect 1273 -710 1277 -707
rect 645 -714 647 -711
rect 786 -714 788 -711
rect 709 -717 711 -714
rect 645 -743 647 -734
rect 850 -717 852 -714
rect 975 -717 990 -713
rect 1114 -714 1116 -711
rect 630 -745 647 -743
rect 630 -747 648 -745
rect 709 -746 711 -737
rect 786 -743 788 -734
rect 986 -720 990 -717
rect 644 -750 648 -747
rect 694 -750 711 -746
rect 771 -745 788 -743
rect 771 -747 789 -745
rect 850 -746 852 -737
rect 1262 -723 1277 -719
rect 1273 -726 1277 -723
rect 986 -743 990 -740
rect 1114 -743 1116 -734
rect 785 -750 789 -747
rect 835 -750 852 -746
rect 1101 -747 1116 -743
rect 1273 -749 1277 -746
rect 724 -762 728 -759
rect 644 -773 648 -770
rect 975 -757 990 -753
rect 865 -762 869 -759
rect 986 -760 990 -757
rect 1103 -760 1107 -757
rect 1154 -760 1158 -757
rect 785 -773 789 -770
rect 724 -785 728 -782
rect 865 -785 869 -782
rect 986 -783 990 -780
rect 1103 -783 1107 -780
rect 1154 -783 1158 -780
rect 711 -789 728 -785
rect 852 -789 869 -785
rect 1090 -787 1107 -783
rect 1141 -787 1158 -783
rect 645 -813 647 -810
rect 701 -813 703 -810
rect 757 -813 759 -810
rect 853 -812 855 -809
rect 909 -812 911 -809
rect 965 -812 967 -809
rect 1021 -812 1023 -809
rect 1145 -812 1147 -809
rect 1201 -812 1203 -809
rect 1257 -812 1259 -809
rect 1313 -812 1315 -809
rect 645 -842 647 -833
rect 701 -842 703 -833
rect 757 -842 759 -833
rect 853 -841 855 -832
rect 909 -841 911 -832
rect 965 -841 967 -832
rect 1021 -841 1023 -832
rect 1145 -841 1147 -832
rect 1201 -841 1203 -832
rect 1257 -841 1259 -832
rect 1313 -841 1315 -832
rect 632 -846 647 -842
rect 688 -846 703 -842
rect 744 -846 759 -842
rect 840 -845 855 -841
rect 896 -845 911 -841
rect 952 -845 967 -841
rect 1008 -845 1023 -841
rect 1132 -845 1147 -841
rect 1188 -845 1203 -841
rect 1244 -845 1259 -841
rect 1300 -845 1315 -841
rect 660 -862 675 -858
rect 868 -861 883 -857
rect 1160 -861 1175 -857
rect 671 -865 675 -862
rect 879 -864 883 -861
rect 1171 -864 1175 -861
rect 671 -888 675 -885
rect 879 -887 883 -884
rect 1171 -887 1175 -884
rect 1427 -890 1429 -887
rect 1483 -890 1485 -887
rect 660 -902 675 -898
rect 868 -901 883 -897
rect 1160 -901 1175 -897
rect 671 -905 675 -902
rect 879 -904 883 -901
rect 1171 -904 1175 -901
rect 1538 -899 1540 -896
rect 1427 -919 1429 -910
rect 1483 -919 1485 -910
rect 1414 -923 1429 -919
rect 1470 -923 1485 -919
rect 671 -928 675 -925
rect 879 -927 883 -924
rect 1171 -927 1175 -924
rect 1538 -928 1540 -919
rect 1523 -930 1540 -928
rect 1523 -932 1541 -930
rect 1537 -935 1541 -932
rect 660 -942 675 -938
rect 868 -941 883 -937
rect 1160 -941 1175 -937
rect 1442 -939 1457 -935
rect 671 -945 675 -942
rect 879 -944 883 -941
rect 1171 -944 1175 -941
rect 1453 -942 1457 -939
rect 1537 -958 1541 -955
rect 671 -968 675 -965
rect 879 -967 883 -964
rect 1171 -967 1175 -964
rect 1453 -965 1457 -962
rect 868 -980 883 -976
rect 1160 -980 1175 -976
rect 1442 -979 1457 -975
rect 879 -983 883 -980
rect 1171 -983 1175 -980
rect 1453 -982 1457 -979
rect 879 -1006 883 -1003
rect 1171 -1006 1175 -1003
rect 1453 -1005 1457 -1002
<< polycontact >>
rect 462 550 466 554
rect 518 550 522 554
rect 637 550 641 554
rect 693 550 697 554
rect 812 550 816 554
rect 868 550 872 554
rect 987 550 991 554
rect 1043 550 1047 554
rect 1165 550 1169 554
rect 1221 550 1225 554
rect 1335 550 1339 554
rect 1391 550 1395 554
rect 1505 550 1509 554
rect 1561 550 1565 554
rect 1675 550 1679 554
rect 1731 550 1735 554
rect 571 541 575 545
rect 746 541 750 545
rect 921 541 925 545
rect 1096 541 1100 545
rect 1274 541 1278 545
rect 1444 541 1448 545
rect 1614 541 1618 545
rect 1784 541 1788 545
rect 490 534 494 538
rect 665 534 669 538
rect 840 534 844 538
rect 1015 534 1019 538
rect 1193 534 1197 538
rect 1363 534 1367 538
rect 1533 534 1537 538
rect 1703 534 1707 538
rect 490 494 494 498
rect 665 494 669 498
rect 840 494 844 498
rect 1015 494 1019 498
rect 1193 494 1197 498
rect 1363 494 1367 498
rect 1533 494 1537 498
rect 1703 494 1707 498
rect 462 399 466 403
rect 518 399 522 403
rect 637 399 641 403
rect 693 399 697 403
rect 812 399 816 403
rect 868 399 872 403
rect 987 399 991 403
rect 1043 399 1047 403
rect 571 390 575 394
rect 746 390 750 394
rect 921 390 925 394
rect 1096 390 1100 394
rect 490 383 494 387
rect 665 383 669 387
rect 840 383 844 387
rect 1015 383 1019 387
rect 490 343 494 347
rect 665 343 669 347
rect 840 343 844 347
rect 1015 343 1019 347
rect 2467 341 2471 345
rect 2530 341 2534 345
rect 2645 341 2649 345
rect 2708 341 2712 345
rect 2800 341 2804 345
rect 2863 341 2867 345
rect 2956 341 2960 345
rect 3019 341 3023 345
rect 2351 305 2355 309
rect 2547 302 2551 306
rect 2725 302 2729 306
rect 2880 302 2884 306
rect 3036 302 3040 306
rect 2531 256 2535 260
rect 2709 256 2713 260
rect 2864 256 2868 260
rect 3020 256 3024 260
rect 1160 239 1164 243
rect 1216 239 1220 243
rect 1335 239 1339 243
rect 1391 239 1395 243
rect 1510 239 1514 243
rect 1566 239 1570 243
rect 1685 239 1689 243
rect 1741 239 1745 243
rect 1269 230 1273 234
rect 1444 230 1448 234
rect 1619 230 1623 234
rect 1794 230 1798 234
rect 616 226 620 230
rect 672 226 676 230
rect 786 226 790 230
rect 842 226 846 230
rect 1188 223 1192 227
rect 725 217 729 221
rect 895 217 899 221
rect 644 210 648 214
rect 814 210 818 214
rect 1363 223 1367 227
rect 1538 223 1542 227
rect 1713 223 1717 227
rect 2548 217 2552 221
rect 2726 217 2730 221
rect 2881 217 2885 221
rect 3037 217 3041 221
rect 1188 183 1192 187
rect 1363 183 1367 187
rect 1538 183 1542 187
rect 1713 183 1717 187
rect 556 170 560 174
rect 644 170 648 174
rect 814 170 818 174
rect 2640 132 2644 136
rect 3162 132 3166 136
rect 2265 128 2269 132
rect 2321 128 2325 132
rect 2447 128 2451 132
rect 2503 128 2507 132
rect 2787 128 2791 132
rect 2843 128 2847 132
rect 2969 128 2973 132
rect 3025 128 3029 132
rect 1007 92 1011 96
rect 2374 119 2378 123
rect 2556 119 2560 123
rect 2896 119 2900 123
rect 3078 119 3082 123
rect 2293 112 2297 116
rect 616 88 620 92
rect 672 88 676 92
rect 786 88 790 92
rect 842 88 846 92
rect 1160 88 1164 92
rect 1216 88 1220 92
rect 1335 88 1339 92
rect 1391 88 1395 92
rect 1510 88 1514 92
rect 1566 88 1570 92
rect 1685 88 1689 92
rect 1741 88 1745 92
rect 2475 112 2479 116
rect 2815 112 2819 116
rect 2640 86 2644 90
rect 2997 112 3001 116
rect 3162 86 3166 90
rect 725 79 729 83
rect 895 79 899 83
rect 1269 79 1273 83
rect 1444 79 1448 83
rect 1619 79 1623 83
rect 1794 79 1798 83
rect 2726 79 2730 83
rect 3248 79 3252 83
rect 644 72 648 76
rect 814 72 818 76
rect 1188 72 1192 76
rect 1007 46 1011 50
rect 1363 72 1367 76
rect 1538 72 1542 76
rect 1713 72 1717 76
rect 2293 72 2297 76
rect 2475 72 2479 76
rect 2815 72 2819 76
rect 2997 72 3001 76
rect 2629 46 2633 50
rect 2680 46 2684 50
rect 3151 46 3155 50
rect 3202 46 3206 50
rect 1093 39 1097 43
rect 556 32 560 36
rect 644 32 648 36
rect 814 32 818 36
rect 1188 32 1192 36
rect 1363 32 1367 36
rect 1538 32 1542 36
rect 1713 32 1717 36
rect 996 6 1000 10
rect 1047 6 1051 10
rect 2322 -10 2326 -6
rect 2385 -10 2389 -6
rect 2633 -7 2637 -3
rect 2696 -7 2700 -3
rect 2844 -10 2848 -6
rect 2907 -10 2911 -6
rect 3155 -7 3159 -3
rect 3218 -7 3222 -3
rect 2402 -49 2406 -45
rect 2713 -46 2717 -42
rect 2924 -49 2928 -45
rect 3235 -46 3239 -42
rect 2322 -92 2326 -88
rect 2633 -89 2637 -85
rect 2386 -95 2390 -91
rect 2697 -92 2701 -88
rect 2844 -92 2848 -88
rect 3155 -89 3159 -85
rect 2908 -95 2912 -91
rect 3219 -92 3223 -88
rect 2403 -134 2407 -130
rect 2714 -131 2718 -127
rect 2925 -134 2929 -130
rect 3236 -131 3240 -127
rect 505 -158 509 -154
rect 561 -158 565 -154
rect 680 -158 684 -154
rect 736 -158 740 -154
rect 855 -158 859 -154
rect 911 -158 915 -154
rect 1030 -158 1034 -154
rect 1086 -158 1090 -154
rect 614 -167 618 -163
rect 789 -167 793 -163
rect 964 -167 968 -163
rect 1139 -167 1143 -163
rect 533 -174 537 -170
rect 708 -174 712 -170
rect 883 -174 887 -170
rect 1058 -174 1062 -170
rect 533 -214 537 -210
rect 708 -214 712 -210
rect 883 -214 887 -210
rect 1058 -214 1062 -210
rect 2640 -254 2644 -250
rect 3162 -254 3166 -250
rect 2265 -258 2269 -254
rect 2321 -258 2325 -254
rect 2447 -258 2451 -254
rect 2503 -258 2507 -254
rect 2787 -258 2791 -254
rect 2843 -258 2847 -254
rect 2969 -258 2973 -254
rect 3025 -258 3029 -254
rect 2374 -267 2378 -263
rect 2556 -267 2560 -263
rect 2896 -267 2900 -263
rect 3078 -267 3082 -263
rect 2293 -274 2297 -270
rect 2475 -274 2479 -270
rect 2815 -274 2819 -270
rect 2640 -300 2644 -296
rect 2997 -274 3001 -270
rect 3162 -300 3166 -296
rect 505 -309 509 -305
rect 561 -309 565 -305
rect 680 -309 684 -305
rect 736 -309 740 -305
rect 855 -309 859 -305
rect 911 -309 915 -305
rect 1030 -309 1034 -305
rect 1086 -309 1090 -305
rect 2726 -307 2730 -303
rect 3248 -307 3252 -303
rect 2293 -314 2297 -310
rect 2475 -314 2479 -310
rect 614 -318 618 -314
rect 789 -318 793 -314
rect 964 -318 968 -314
rect 1139 -318 1143 -314
rect 533 -325 537 -321
rect 708 -325 712 -321
rect 883 -325 887 -321
rect 1058 -325 1062 -321
rect 2815 -314 2819 -310
rect 2997 -314 3001 -310
rect 2629 -340 2633 -336
rect 2680 -340 2684 -336
rect 3151 -340 3155 -336
rect 3202 -340 3206 -336
rect 533 -365 537 -361
rect 708 -365 712 -361
rect 883 -365 887 -361
rect 1058 -365 1062 -361
rect 2322 -396 2326 -392
rect 2385 -396 2389 -392
rect 2633 -393 2637 -389
rect 2696 -393 2700 -389
rect 2844 -396 2848 -392
rect 2907 -396 2911 -392
rect 3155 -393 3159 -389
rect 3218 -393 3222 -389
rect 2402 -435 2406 -431
rect 2713 -432 2717 -428
rect 2924 -435 2928 -431
rect 3235 -432 3239 -428
rect 2322 -478 2326 -474
rect 2633 -475 2637 -471
rect 626 -484 630 -480
rect 689 -484 693 -480
rect 767 -484 771 -480
rect 830 -484 834 -480
rect 913 -484 917 -480
rect 969 -484 973 -480
rect 1025 -484 1029 -480
rect 1081 -484 1085 -480
rect 2386 -481 2390 -477
rect 2697 -478 2701 -474
rect 2844 -478 2848 -474
rect 3155 -475 3159 -471
rect 1131 -493 1135 -489
rect 941 -500 945 -496
rect 706 -523 710 -519
rect 847 -523 851 -519
rect 2908 -481 2912 -477
rect 3219 -478 3223 -474
rect 2403 -520 2407 -516
rect 2714 -517 2718 -513
rect 2925 -520 2929 -516
rect 3236 -517 3240 -513
rect 626 -566 630 -562
rect 941 -540 945 -536
rect 690 -569 694 -565
rect 767 -566 771 -562
rect 1230 -549 1234 -545
rect 1286 -549 1290 -545
rect 1342 -549 1346 -545
rect 1398 -549 1402 -545
rect 1453 -549 1457 -545
rect 831 -569 835 -565
rect 1258 -565 1262 -561
rect 941 -580 945 -576
rect 707 -608 711 -604
rect 848 -608 852 -604
rect 1258 -605 1262 -601
rect 941 -619 945 -615
rect 1592 -620 1596 -616
rect 1648 -620 1652 -616
rect 1762 -620 1766 -616
rect 1818 -620 1822 -616
rect 1932 -620 1936 -616
rect 1988 -620 1992 -616
rect 2102 -620 2106 -616
rect 2158 -620 2162 -616
rect 1701 -629 1705 -625
rect 1871 -629 1875 -625
rect 2041 -629 2045 -625
rect 2211 -629 2215 -625
rect 1620 -636 1624 -632
rect 1258 -645 1262 -641
rect 626 -665 630 -661
rect 689 -665 693 -661
rect 767 -665 771 -661
rect 830 -665 834 -661
rect 1790 -636 1794 -632
rect 1960 -636 1964 -632
rect 2130 -636 2134 -632
rect 1620 -676 1624 -672
rect 1790 -676 1794 -672
rect 1960 -676 1964 -672
rect 2130 -676 2134 -672
rect 1258 -684 1262 -680
rect 706 -704 710 -700
rect 847 -704 851 -700
rect 943 -701 947 -697
rect 999 -701 1003 -697
rect 1097 -701 1101 -697
rect 971 -717 975 -713
rect 626 -747 630 -743
rect 690 -750 694 -746
rect 767 -747 771 -743
rect 1258 -723 1262 -719
rect 831 -750 835 -746
rect 1097 -747 1101 -743
rect 971 -757 975 -753
rect 707 -789 711 -785
rect 848 -789 852 -785
rect 1086 -787 1090 -783
rect 1137 -787 1141 -783
rect 628 -846 632 -842
rect 684 -846 688 -842
rect 740 -846 744 -842
rect 836 -845 840 -841
rect 892 -845 896 -841
rect 948 -845 952 -841
rect 1004 -845 1008 -841
rect 1128 -845 1132 -841
rect 1184 -845 1188 -841
rect 1240 -845 1244 -841
rect 1296 -845 1300 -841
rect 656 -862 660 -858
rect 864 -861 868 -857
rect 1156 -861 1160 -857
rect 656 -902 660 -898
rect 864 -901 868 -897
rect 1156 -901 1160 -897
rect 1410 -923 1414 -919
rect 1466 -923 1470 -919
rect 1519 -932 1523 -928
rect 656 -942 660 -938
rect 864 -941 868 -937
rect 1156 -941 1160 -937
rect 1438 -939 1442 -935
rect 864 -980 868 -976
rect 1156 -980 1160 -976
rect 1438 -979 1442 -975
<< metal1 >>
rect 447 597 622 602
rect 627 597 797 602
rect 802 597 972 602
rect 447 554 452 597
rect 466 589 550 593
rect 554 589 573 593
rect 577 589 605 593
rect 609 589 637 593
rect 641 589 725 593
rect 729 589 748 593
rect 752 589 780 593
rect 784 589 812 593
rect 816 589 900 593
rect 904 589 923 593
rect 927 589 955 593
rect 959 589 987 593
rect 991 589 1075 593
rect 1079 589 1098 593
rect 1102 589 1130 593
rect 1169 589 1253 593
rect 1257 589 1276 593
rect 1280 589 1308 593
rect 1312 589 1335 593
rect 1339 589 1423 593
rect 1427 589 1446 593
rect 1450 589 1478 593
rect 1482 589 1505 593
rect 1509 589 1593 593
rect 1597 589 1616 593
rect 1620 589 1648 593
rect 1652 589 1675 593
rect 1679 589 1763 593
rect 1767 589 1786 593
rect 1790 589 1818 593
rect 468 583 478 589
rect 524 583 534 589
rect 447 550 462 554
rect 447 538 452 550
rect 482 545 492 563
rect 503 550 518 554
rect 538 545 548 563
rect 579 574 589 589
rect 643 583 653 589
rect 699 583 709 589
rect 594 545 603 554
rect 627 550 637 554
rect 462 541 571 545
rect 594 541 617 545
rect 447 534 490 538
rect 447 403 452 534
rect 510 531 520 541
rect 594 538 603 541
rect 622 538 627 550
rect 657 545 667 563
rect 678 550 693 554
rect 713 545 723 563
rect 754 574 764 589
rect 818 583 828 589
rect 874 583 884 589
rect 769 545 778 554
rect 802 550 812 554
rect 637 541 746 545
rect 769 541 792 545
rect 622 534 665 538
rect 685 531 695 541
rect 769 538 778 541
rect 797 538 802 550
rect 832 545 842 563
rect 853 550 868 554
rect 888 545 898 563
rect 929 574 939 589
rect 993 583 1003 589
rect 1049 583 1059 589
rect 944 545 953 554
rect 977 550 987 554
rect 812 541 921 545
rect 944 541 967 545
rect 494 505 504 511
rect 494 501 520 505
rect 475 494 490 498
rect 510 491 520 501
rect 494 465 504 471
rect 578 465 588 518
rect 797 534 840 538
rect 860 531 870 541
rect 944 538 953 541
rect 972 538 977 550
rect 1007 545 1017 563
rect 1028 550 1043 554
rect 1063 545 1073 563
rect 1104 574 1114 589
rect 1171 583 1181 589
rect 1227 583 1237 589
rect 1119 545 1128 554
rect 1150 550 1165 554
rect 1185 545 1195 563
rect 1206 550 1221 554
rect 1241 545 1251 563
rect 1282 574 1292 589
rect 1341 583 1351 589
rect 1397 583 1407 589
rect 1297 545 1306 554
rect 1320 550 1335 554
rect 1355 545 1365 563
rect 1376 550 1391 554
rect 1411 545 1421 563
rect 1452 574 1462 589
rect 1511 583 1521 589
rect 1567 583 1577 589
rect 1467 545 1476 554
rect 1490 550 1505 554
rect 1525 545 1535 563
rect 1546 550 1561 554
rect 1581 545 1591 563
rect 1622 574 1632 589
rect 1681 583 1691 589
rect 1737 583 1747 589
rect 1637 545 1646 554
rect 1660 550 1675 554
rect 1695 545 1705 563
rect 1716 550 1731 554
rect 1751 545 1761 563
rect 1792 574 1802 589
rect 1807 545 1816 554
rect 987 541 1096 545
rect 1119 541 1142 545
rect 1165 541 1274 545
rect 1297 541 1320 545
rect 1335 541 1444 545
rect 1467 541 1490 545
rect 1505 541 1614 545
rect 1637 541 1660 545
rect 1675 541 1784 545
rect 1807 541 1830 545
rect 669 505 679 511
rect 669 501 695 505
rect 650 494 665 498
rect 685 491 695 501
rect 669 465 679 471
rect 753 465 763 518
rect 972 534 1015 538
rect 1035 531 1045 541
rect 1119 538 1128 541
rect 844 505 854 511
rect 844 501 870 505
rect 825 494 840 498
rect 860 491 870 501
rect 844 465 854 471
rect 928 465 938 518
rect 1178 534 1193 538
rect 1213 531 1223 541
rect 1297 538 1306 541
rect 1019 505 1029 511
rect 1019 501 1045 505
rect 1000 494 1015 498
rect 1035 491 1045 501
rect 1019 465 1029 471
rect 1103 465 1113 518
rect 1348 534 1363 538
rect 1383 531 1393 541
rect 1467 538 1476 541
rect 1197 505 1207 511
rect 1197 501 1223 505
rect 1178 494 1193 498
rect 1213 491 1223 501
rect 1197 465 1207 471
rect 1281 465 1291 518
rect 1518 534 1533 538
rect 1553 531 1563 541
rect 1637 538 1646 541
rect 1367 505 1377 511
rect 1367 501 1393 505
rect 1348 494 1363 498
rect 1383 491 1393 501
rect 1367 465 1377 471
rect 1451 465 1461 518
rect 1688 534 1703 538
rect 1723 531 1733 541
rect 1807 538 1816 541
rect 1537 505 1547 511
rect 1537 501 1563 505
rect 1518 494 1533 498
rect 1553 491 1563 501
rect 1537 465 1547 471
rect 1621 465 1631 518
rect 1707 505 1717 511
rect 1707 501 1733 505
rect 1688 494 1703 498
rect 1723 491 1733 501
rect 1707 465 1717 471
rect 1791 465 1801 518
rect 466 461 550 465
rect 554 461 573 465
rect 577 461 605 465
rect 609 461 637 465
rect 641 461 725 465
rect 729 461 748 465
rect 752 461 780 465
rect 784 461 812 465
rect 816 461 900 465
rect 904 461 923 465
rect 927 461 955 465
rect 959 461 987 465
rect 991 461 1075 465
rect 1079 461 1098 465
rect 1102 461 1130 465
rect 1169 461 1253 465
rect 1257 461 1276 465
rect 1280 461 1308 465
rect 1312 461 1335 465
rect 1339 461 1423 465
rect 1427 461 1446 465
rect 1450 461 1478 465
rect 1482 461 1505 465
rect 1509 461 1593 465
rect 1597 461 1616 465
rect 1620 461 1648 465
rect 1652 461 1675 465
rect 1679 461 1763 465
rect 1767 461 1786 465
rect 1790 461 1818 465
rect 466 438 550 442
rect 554 438 573 442
rect 577 438 605 442
rect 609 438 637 442
rect 641 438 725 442
rect 729 438 748 442
rect 752 438 780 442
rect 784 438 812 442
rect 816 438 900 442
rect 904 438 923 442
rect 927 438 955 442
rect 959 438 987 442
rect 991 438 1075 442
rect 1079 438 1098 442
rect 1102 438 1130 442
rect 468 432 478 438
rect 524 432 534 438
rect 447 399 462 403
rect 447 387 452 399
rect 482 394 492 412
rect 503 399 518 403
rect 538 394 548 412
rect 579 423 589 438
rect 643 432 653 438
rect 699 432 709 438
rect 594 394 603 403
rect 622 399 637 403
rect 462 390 571 394
rect 594 390 617 394
rect 447 383 490 387
rect 447 296 452 383
rect 510 380 520 390
rect 594 387 603 390
rect 622 388 627 399
rect 657 394 667 412
rect 678 399 693 403
rect 713 394 723 412
rect 754 423 764 438
rect 818 432 828 438
rect 874 432 884 438
rect 769 394 778 403
rect 797 399 812 403
rect 637 390 746 394
rect 769 390 792 394
rect 627 383 665 387
rect 685 380 695 390
rect 769 387 778 390
rect 797 388 802 399
rect 832 394 842 412
rect 853 399 868 403
rect 888 394 898 412
rect 929 423 939 438
rect 993 432 1003 438
rect 1049 432 1059 438
rect 944 394 953 403
rect 972 399 987 403
rect 812 390 921 394
rect 944 390 967 394
rect 494 354 504 360
rect 494 350 520 354
rect 475 343 490 347
rect 510 340 520 350
rect 494 314 504 320
rect 578 314 588 367
rect 802 383 840 387
rect 860 380 870 390
rect 944 387 953 390
rect 972 388 977 399
rect 1007 394 1017 412
rect 1028 399 1043 403
rect 1063 394 1073 412
rect 1104 423 1114 438
rect 1119 394 1128 403
rect 987 390 1096 394
rect 1119 390 1142 394
rect 669 354 679 360
rect 669 350 695 354
rect 650 343 665 347
rect 685 340 695 350
rect 669 314 679 320
rect 753 314 763 367
rect 977 383 1015 387
rect 1035 380 1045 390
rect 1119 387 1128 390
rect 844 354 854 360
rect 844 350 870 354
rect 825 343 840 347
rect 860 340 870 350
rect 844 314 854 320
rect 928 314 938 367
rect 2473 380 2501 384
rect 2532 380 2579 384
rect 2651 380 2679 384
rect 2710 380 2757 384
rect 2806 380 2834 384
rect 2865 380 2912 384
rect 2962 380 2990 384
rect 3021 380 3068 384
rect 2475 374 2485 380
rect 2538 374 2548 380
rect 1019 354 1029 360
rect 1019 350 1045 354
rect 1000 343 1015 347
rect 1035 340 1045 350
rect 1019 314 1029 320
rect 1103 314 1113 367
rect 2357 344 2385 348
rect 2490 345 2499 354
rect 2359 338 2369 344
rect 2453 341 2467 345
rect 2490 341 2513 345
rect 2517 341 2530 345
rect 2490 338 2499 341
rect 466 310 550 314
rect 554 310 573 314
rect 577 310 605 314
rect 609 310 637 314
rect 641 310 725 314
rect 729 310 748 314
rect 752 310 780 314
rect 784 310 812 314
rect 816 310 900 314
rect 904 310 923 314
rect 927 310 955 314
rect 959 310 987 314
rect 991 310 1075 314
rect 1079 310 1098 314
rect 1102 310 1130 314
rect 1134 310 1142 314
rect 2374 309 2383 318
rect 2553 329 2562 354
rect 2569 329 2579 380
rect 2653 374 2663 380
rect 2716 374 2726 380
rect 2668 345 2677 354
rect 2631 341 2645 345
rect 2668 341 2691 345
rect 2695 341 2708 345
rect 2668 338 2677 341
rect 2474 312 2484 318
rect 1145 305 1320 309
rect 447 291 622 296
rect 627 291 766 296
rect 771 291 797 296
rect 802 291 972 296
rect 490 276 946 281
rect 490 -106 495 276
rect 526 265 558 269
rect 562 265 590 269
rect 594 265 616 269
rect 620 265 704 269
rect 708 265 727 269
rect 731 265 759 269
rect 763 265 786 269
rect 790 265 874 269
rect 878 265 897 269
rect 901 265 929 269
rect 526 131 530 265
rect 564 203 574 265
rect 622 259 632 265
rect 678 259 688 265
rect 601 226 616 230
rect 636 221 646 239
rect 657 226 672 230
rect 692 221 702 239
rect 733 250 743 265
rect 792 259 802 265
rect 848 259 858 265
rect 748 221 757 230
rect 771 226 786 230
rect 616 217 725 221
rect 748 217 766 221
rect 806 221 816 239
rect 827 226 842 230
rect 862 221 872 239
rect 903 250 913 265
rect 918 221 927 230
rect 941 221 946 276
rect 786 217 895 221
rect 918 217 946 221
rect 1145 243 1149 305
rect 1325 305 1495 309
rect 1500 305 1670 309
rect 2337 305 2351 309
rect 2374 305 2397 309
rect 2473 308 2501 312
rect 2731 329 2740 354
rect 2747 329 2757 380
rect 2808 374 2818 380
rect 2871 374 2881 380
rect 2823 345 2832 354
rect 2786 341 2800 345
rect 2823 341 2846 345
rect 2850 341 2863 345
rect 2823 338 2832 341
rect 2652 312 2662 318
rect 2651 308 2679 312
rect 2886 329 2895 354
rect 2902 329 2912 380
rect 2964 374 2974 380
rect 3027 374 3037 380
rect 2979 345 2988 354
rect 2942 341 2956 345
rect 2979 341 3002 345
rect 3006 341 3019 345
rect 2979 338 2988 341
rect 2807 312 2817 318
rect 2806 308 2834 312
rect 3042 329 3051 354
rect 3058 329 3068 380
rect 2963 312 2973 318
rect 2962 308 2990 312
rect 2374 302 2383 305
rect 2533 302 2547 306
rect 2711 302 2725 306
rect 2866 302 2880 306
rect 3022 302 3036 306
rect 2533 295 2579 299
rect 2711 295 2757 299
rect 2866 295 2912 299
rect 3022 295 3068 299
rect 2539 289 2549 295
rect 1164 278 1248 282
rect 1252 278 1271 282
rect 1275 278 1303 282
rect 1307 278 1335 282
rect 1339 278 1423 282
rect 1427 278 1446 282
rect 1450 278 1478 282
rect 1482 278 1510 282
rect 1514 278 1598 282
rect 1602 278 1621 282
rect 1625 278 1653 282
rect 1657 278 1685 282
rect 1689 278 1773 282
rect 1777 278 1796 282
rect 1800 278 1828 282
rect 1166 272 1176 278
rect 1222 272 1232 278
rect 1145 239 1160 243
rect 1145 227 1149 239
rect 1180 234 1190 252
rect 1201 239 1216 243
rect 1236 234 1246 252
rect 1277 263 1287 278
rect 1341 272 1351 278
rect 1397 272 1407 278
rect 1292 234 1301 243
rect 1325 239 1335 243
rect 1160 230 1269 234
rect 1292 230 1315 234
rect 1145 223 1188 227
rect 629 210 644 214
rect 664 207 674 217
rect 748 214 757 217
rect 579 174 588 183
rect 799 210 814 214
rect 834 207 844 217
rect 918 214 927 217
rect 648 181 658 187
rect 648 177 674 181
rect 542 170 556 174
rect 579 170 602 174
rect 629 170 644 174
rect 579 167 588 170
rect 664 167 674 177
rect 563 141 573 147
rect 648 141 658 147
rect 732 141 742 194
rect 818 181 828 187
rect 818 177 844 181
rect 799 170 814 174
rect 834 167 844 177
rect 818 141 828 147
rect 902 141 912 194
rect 562 137 590 141
rect 594 137 616 141
rect 620 137 704 141
rect 708 137 727 141
rect 731 137 759 141
rect 763 137 786 141
rect 790 137 874 141
rect 878 137 897 141
rect 901 137 929 141
rect 933 137 965 141
rect 526 127 558 131
rect 562 127 590 131
rect 594 127 616 131
rect 620 127 704 131
rect 708 127 727 131
rect 731 127 759 131
rect 763 127 786 131
rect 790 127 874 131
rect 878 127 897 131
rect 901 127 929 131
rect 564 65 574 127
rect 622 121 632 127
rect 678 121 688 127
rect 601 88 616 92
rect 636 83 646 101
rect 657 88 672 92
rect 692 83 702 101
rect 733 112 743 127
rect 792 121 802 127
rect 848 121 858 127
rect 748 83 757 92
rect 771 88 786 92
rect 616 79 725 83
rect 748 79 767 83
rect 806 83 816 101
rect 827 88 842 92
rect 862 83 872 101
rect 903 112 913 127
rect 918 83 927 92
rect 786 79 895 83
rect 918 79 937 83
rect 629 72 644 76
rect 664 69 674 79
rect 748 76 757 79
rect 579 36 588 45
rect 799 72 814 76
rect 834 69 844 79
rect 918 76 927 79
rect 648 43 658 49
rect 648 39 674 43
rect 543 32 556 36
rect 579 32 602 36
rect 629 32 644 36
rect 579 29 588 32
rect 664 29 674 39
rect 563 3 573 9
rect 648 3 658 9
rect 732 3 742 56
rect 818 43 828 49
rect 818 39 844 43
rect 799 32 814 36
rect 834 29 844 39
rect 818 3 828 9
rect 902 3 912 56
rect 961 3 965 137
rect 982 131 1007 135
rect 1011 131 1039 135
rect 1043 131 1095 135
rect 1099 131 1127 135
rect 1013 125 1023 131
rect 997 92 1007 96
rect 1027 89 1037 105
rect 1007 85 1043 89
rect 1013 79 1023 85
rect 997 46 1007 50
rect 1027 43 1037 59
rect 1101 72 1111 131
rect 1145 92 1149 223
rect 1208 220 1218 230
rect 1292 227 1301 230
rect 1320 227 1325 239
rect 1355 234 1365 252
rect 1376 239 1391 243
rect 1411 234 1421 252
rect 1452 263 1462 278
rect 1516 272 1526 278
rect 1572 272 1582 278
rect 1467 234 1476 243
rect 1500 239 1510 243
rect 1335 230 1444 234
rect 1467 230 1490 234
rect 1320 223 1363 227
rect 1383 220 1393 230
rect 1467 227 1476 230
rect 1495 227 1500 239
rect 1530 234 1540 252
rect 1551 239 1566 243
rect 1586 234 1596 252
rect 1627 263 1637 278
rect 1691 272 1701 278
rect 1747 272 1757 278
rect 1642 234 1651 243
rect 1675 239 1685 243
rect 1510 230 1619 234
rect 1642 230 1665 234
rect 1192 194 1202 200
rect 1192 190 1218 194
rect 1173 183 1188 187
rect 1208 180 1218 190
rect 1192 154 1202 160
rect 1276 154 1286 207
rect 1495 223 1538 227
rect 1558 220 1568 230
rect 1642 227 1651 230
rect 1670 227 1675 239
rect 1705 234 1715 252
rect 1726 239 1741 243
rect 1761 234 1771 252
rect 1802 263 1812 278
rect 2358 276 2368 282
rect 2357 272 2385 276
rect 2517 256 2531 260
rect 1817 234 1826 243
rect 2554 244 2563 269
rect 2570 244 2579 295
rect 2717 289 2727 295
rect 2695 256 2709 260
rect 1685 230 1794 234
rect 1817 230 1840 234
rect 1367 194 1377 200
rect 1367 190 1393 194
rect 1348 183 1363 187
rect 1383 180 1393 190
rect 1367 154 1377 160
rect 1451 154 1461 207
rect 1670 223 1713 227
rect 1733 220 1743 230
rect 1817 227 1826 230
rect 1542 194 1552 200
rect 1542 190 1568 194
rect 1523 183 1538 187
rect 1558 180 1568 190
rect 1542 154 1552 160
rect 1626 154 1636 207
rect 2732 244 2741 269
rect 2748 244 2757 295
rect 2872 289 2882 295
rect 2850 256 2864 260
rect 2887 244 2896 269
rect 2903 244 2912 295
rect 3028 289 3038 295
rect 3006 256 3020 260
rect 3043 244 3052 269
rect 3059 244 3068 295
rect 2534 217 2548 221
rect 2712 217 2726 221
rect 2867 217 2881 221
rect 3023 217 3037 221
rect 1717 194 1727 200
rect 1717 190 1743 194
rect 1698 183 1713 187
rect 1733 180 1743 190
rect 1717 154 1727 160
rect 1801 154 1811 207
rect 2269 171 2353 175
rect 2357 171 2376 175
rect 2380 171 2408 175
rect 2412 171 2447 175
rect 2451 171 2535 175
rect 2539 171 2558 175
rect 2562 171 2590 175
rect 2594 171 2640 175
rect 2644 171 2672 175
rect 2676 171 2728 175
rect 2732 171 2760 175
rect 2764 171 2787 175
rect 2791 171 2875 175
rect 2879 171 2898 175
rect 2902 171 2930 175
rect 2934 171 2969 175
rect 2973 171 3057 175
rect 3061 171 3080 175
rect 3084 171 3112 175
rect 3116 171 3162 175
rect 3166 171 3194 175
rect 3198 171 3250 175
rect 3254 171 3282 175
rect 2271 161 2281 171
rect 2327 161 2337 171
rect 1164 150 1248 154
rect 1252 150 1271 154
rect 1275 150 1303 154
rect 1307 150 1335 154
rect 1339 150 1423 154
rect 1427 150 1446 154
rect 1450 150 1478 154
rect 1482 150 1510 154
rect 1514 150 1598 154
rect 1602 150 1621 154
rect 1625 150 1653 154
rect 1657 150 1685 154
rect 1689 150 1773 154
rect 1777 150 1796 154
rect 1800 150 1828 154
rect 1164 127 1248 131
rect 1252 127 1271 131
rect 1275 127 1303 131
rect 1307 127 1335 131
rect 1339 127 1423 131
rect 1427 127 1446 131
rect 1450 127 1478 131
rect 1482 127 1510 131
rect 1514 127 1598 131
rect 1602 127 1621 131
rect 1625 127 1653 131
rect 1657 127 1685 131
rect 1689 127 1773 131
rect 1777 127 1796 131
rect 1800 127 1828 131
rect 2250 128 2265 132
rect 1166 121 1176 127
rect 1222 121 1232 127
rect 1145 88 1160 92
rect 1145 76 1149 88
rect 1180 83 1190 101
rect 1201 88 1216 92
rect 1236 83 1246 101
rect 1277 112 1287 127
rect 1341 121 1351 127
rect 1397 121 1407 127
rect 1292 83 1301 92
rect 1320 88 1335 92
rect 1160 79 1269 83
rect 1292 79 1315 83
rect 1145 72 1188 76
rect 1116 43 1125 52
rect 1173 43 1177 72
rect 1208 69 1218 79
rect 1292 76 1301 79
rect 1320 77 1325 88
rect 1355 83 1365 101
rect 1376 88 1391 92
rect 1411 83 1421 101
rect 1452 112 1462 127
rect 1516 121 1526 127
rect 1572 121 1582 127
rect 1467 83 1476 92
rect 1495 88 1510 92
rect 1335 79 1444 83
rect 1467 79 1490 83
rect 982 39 1093 43
rect 1116 39 1177 43
rect 1325 72 1363 76
rect 1383 69 1393 79
rect 1467 76 1476 79
rect 1495 77 1500 88
rect 1530 83 1540 101
rect 1551 88 1566 92
rect 1586 83 1596 101
rect 1627 112 1637 127
rect 1691 121 1701 127
rect 1747 121 1757 127
rect 1642 83 1651 92
rect 1670 88 1685 92
rect 1510 79 1619 83
rect 1642 79 1665 83
rect 1192 43 1202 49
rect 1192 39 1218 43
rect 1002 33 1012 39
rect 1053 33 1063 39
rect 1116 36 1125 39
rect 986 6 996 10
rect 1018 3 1028 13
rect 1038 6 1047 10
rect 1069 3 1079 13
rect 1100 3 1110 16
rect 562 -1 590 3
rect 594 -1 616 3
rect 620 -1 704 3
rect 708 -1 727 3
rect 731 -1 759 3
rect 763 -1 786 3
rect 790 -1 874 3
rect 878 -1 897 3
rect 901 -1 929 3
rect 933 -1 965 3
rect 986 -1 1075 3
rect 1079 -1 1095 3
rect 1099 -1 1127 3
rect 1145 -23 1149 39
rect 1173 32 1188 36
rect 1208 29 1218 39
rect 1192 3 1202 9
rect 1276 3 1286 56
rect 1500 72 1538 76
rect 1558 69 1568 79
rect 1642 76 1651 79
rect 1670 77 1675 88
rect 1705 83 1715 101
rect 1726 88 1741 92
rect 1761 83 1771 101
rect 1802 112 1812 127
rect 2285 123 2295 141
rect 2306 128 2321 132
rect 2341 123 2351 141
rect 2382 152 2392 171
rect 2453 161 2463 171
rect 2509 161 2519 171
rect 2397 123 2406 132
rect 2432 128 2447 132
rect 2467 123 2477 141
rect 2488 128 2503 132
rect 2523 123 2533 141
rect 2564 152 2574 171
rect 2646 165 2656 171
rect 2626 132 2640 136
rect 2579 123 2588 132
rect 2660 129 2670 145
rect 2640 125 2676 129
rect 2265 119 2374 123
rect 2397 119 2420 123
rect 2447 119 2556 123
rect 2579 119 2602 123
rect 2646 119 2656 125
rect 2278 112 2293 116
rect 2313 109 2323 119
rect 2397 116 2406 119
rect 1817 83 1826 92
rect 2460 112 2475 116
rect 2495 109 2505 119
rect 2579 116 2588 119
rect 2297 83 2307 89
rect 1685 79 1794 83
rect 1817 79 1840 83
rect 2297 79 2323 83
rect 1367 43 1377 49
rect 1367 39 1393 43
rect 1348 32 1363 36
rect 1383 29 1393 39
rect 1367 3 1377 9
rect 1451 3 1461 56
rect 1675 72 1713 76
rect 1733 69 1743 79
rect 1817 76 1826 79
rect 1542 43 1552 49
rect 1542 39 1568 43
rect 1523 32 1538 36
rect 1558 29 1568 39
rect 1542 3 1552 9
rect 1626 3 1636 56
rect 2278 72 2293 76
rect 2313 69 2323 79
rect 1717 43 1727 49
rect 1717 39 1743 43
rect 1698 32 1713 36
rect 1733 29 1743 39
rect 1717 3 1727 9
rect 1801 3 1811 56
rect 2297 43 2307 49
rect 2381 43 2391 96
rect 2479 83 2489 89
rect 2479 79 2505 83
rect 2460 72 2475 76
rect 2495 69 2505 79
rect 2479 43 2489 49
rect 2563 43 2573 96
rect 2626 86 2640 90
rect 2660 83 2670 99
rect 2734 112 2744 171
rect 2793 161 2803 171
rect 2849 161 2859 171
rect 2772 128 2787 132
rect 2807 123 2817 141
rect 2828 128 2843 132
rect 2863 123 2873 141
rect 2904 152 2914 171
rect 2975 161 2985 171
rect 3031 161 3041 171
rect 2919 123 2928 132
rect 2954 128 2969 132
rect 2989 123 2999 141
rect 3010 128 3025 132
rect 3045 123 3055 141
rect 3086 152 3096 171
rect 3168 165 3178 171
rect 3148 132 3162 136
rect 3101 123 3110 132
rect 3182 129 3192 145
rect 3162 125 3198 129
rect 2787 119 2896 123
rect 2919 119 2942 123
rect 2969 119 3078 123
rect 3101 119 3124 123
rect 3168 119 3178 125
rect 2800 112 2815 116
rect 2835 109 2845 119
rect 2919 116 2928 119
rect 2749 83 2758 92
rect 2982 112 2997 116
rect 3017 109 3027 119
rect 3101 116 3110 119
rect 2819 83 2829 89
rect 2615 79 2726 83
rect 2749 79 2772 83
rect 2819 79 2845 83
rect 2635 73 2645 79
rect 2686 73 2696 79
rect 2749 76 2758 79
rect 2615 46 2629 50
rect 2651 43 2661 53
rect 2666 46 2680 50
rect 2702 43 2712 53
rect 2800 72 2815 76
rect 2835 69 2845 79
rect 2733 43 2743 56
rect 2819 43 2829 49
rect 2903 43 2913 96
rect 3001 83 3011 89
rect 3001 79 3027 83
rect 2982 72 2997 76
rect 3017 69 3027 79
rect 3001 43 3011 49
rect 3085 43 3095 96
rect 3148 86 3162 90
rect 3182 83 3192 99
rect 3256 112 3266 171
rect 3271 83 3280 92
rect 3137 79 3248 83
rect 3271 79 3294 83
rect 3157 73 3167 79
rect 3208 73 3218 79
rect 3271 76 3280 79
rect 3137 46 3151 50
rect 3173 43 3183 53
rect 3188 46 3202 50
rect 3224 43 3234 53
rect 3255 43 3265 56
rect 2269 39 2353 43
rect 2357 39 2376 43
rect 2380 39 2408 43
rect 2412 39 2447 43
rect 2451 39 2535 43
rect 2539 39 2558 43
rect 2562 39 2590 43
rect 2594 39 2615 43
rect 2619 39 2708 43
rect 2712 39 2728 43
rect 2732 39 2760 43
rect 2764 39 2787 43
rect 2791 39 2875 43
rect 2879 39 2898 43
rect 2902 39 2930 43
rect 2934 39 2969 43
rect 2973 39 3057 43
rect 3061 39 3080 43
rect 3084 39 3112 43
rect 3116 39 3137 43
rect 3141 39 3230 43
rect 3234 39 3250 43
rect 3254 39 3282 43
rect 2328 29 2356 33
rect 2387 29 2434 33
rect 2639 32 2667 36
rect 2698 32 2745 36
rect 2330 23 2340 29
rect 2393 23 2403 29
rect 1164 -1 1248 3
rect 1252 -1 1271 3
rect 1275 -1 1303 3
rect 1307 -1 1335 3
rect 1339 -1 1423 3
rect 1427 -1 1446 3
rect 1450 -1 1478 3
rect 1482 -1 1510 3
rect 1514 -1 1598 3
rect 1602 -1 1621 3
rect 1625 -1 1653 3
rect 1657 -1 1685 3
rect 1689 -1 1773 3
rect 1777 -1 1796 3
rect 1800 -1 1828 3
rect 1832 -1 1840 3
rect 2345 -6 2354 3
rect 2308 -10 2322 -6
rect 2345 -10 2368 -6
rect 2372 -10 2385 -6
rect 2345 -13 2354 -10
rect 1145 -28 1320 -23
rect 1325 -28 1495 -23
rect 1500 -28 1670 -23
rect 2408 -22 2417 3
rect 2424 -22 2434 29
rect 2641 26 2651 32
rect 2704 26 2714 32
rect 2656 -3 2665 6
rect 2619 -7 2633 -3
rect 2656 -7 2679 -3
rect 2683 -7 2696 -3
rect 2656 -10 2665 -7
rect 2329 -39 2339 -33
rect 2328 -43 2356 -39
rect 2719 -19 2728 6
rect 2735 -19 2745 32
rect 2850 29 2878 33
rect 2909 29 2956 33
rect 3161 32 3189 36
rect 3220 32 3267 36
rect 2852 23 2862 29
rect 2915 23 2925 29
rect 2867 -6 2876 3
rect 2830 -10 2844 -6
rect 2867 -10 2890 -6
rect 2894 -10 2907 -6
rect 2867 -13 2876 -10
rect 2640 -36 2650 -30
rect 2639 -40 2667 -36
rect 2930 -22 2939 3
rect 2946 -22 2956 29
rect 3163 26 3173 32
rect 3226 26 3236 32
rect 3178 -3 3187 6
rect 3141 -7 3155 -3
rect 3178 -7 3201 -3
rect 3205 -7 3218 -3
rect 3178 -10 3187 -7
rect 2851 -39 2861 -33
rect 2388 -49 2402 -45
rect 2699 -46 2713 -42
rect 2850 -43 2878 -39
rect 3241 -19 3250 6
rect 3257 -19 3267 32
rect 3162 -36 3172 -30
rect 3161 -40 3189 -36
rect 2328 -53 2356 -49
rect 2639 -50 2667 -46
rect 2910 -49 2924 -45
rect 3221 -46 3235 -42
rect 2330 -59 2340 -53
rect 2388 -56 2434 -52
rect 2345 -88 2354 -79
rect 2394 -62 2404 -56
rect 2308 -92 2322 -88
rect 2345 -92 2368 -88
rect 2345 -95 2354 -92
rect 2372 -95 2386 -91
rect 490 -111 1020 -106
rect 490 -154 495 -111
rect 2409 -107 2418 -82
rect 2425 -107 2434 -56
rect 2641 -56 2651 -50
rect 2699 -53 2745 -49
rect 2850 -53 2878 -49
rect 3161 -50 3189 -46
rect 2656 -85 2665 -76
rect 2705 -59 2715 -53
rect 2619 -89 2633 -85
rect 2656 -89 2679 -85
rect 2656 -92 2665 -89
rect 2683 -92 2697 -88
rect 509 -119 593 -115
rect 597 -119 616 -115
rect 620 -119 648 -115
rect 652 -119 680 -115
rect 684 -119 768 -115
rect 772 -119 791 -115
rect 795 -119 823 -115
rect 827 -119 855 -115
rect 859 -119 943 -115
rect 947 -119 966 -115
rect 970 -119 998 -115
rect 1002 -119 1030 -115
rect 1034 -119 1118 -115
rect 1122 -119 1141 -115
rect 1145 -119 1173 -115
rect 511 -125 521 -119
rect 567 -125 577 -119
rect 490 -158 505 -154
rect 490 -170 495 -158
rect 525 -163 535 -145
rect 546 -158 561 -154
rect 581 -163 591 -145
rect 622 -134 632 -119
rect 686 -125 696 -119
rect 742 -125 752 -119
rect 637 -163 646 -154
rect 665 -158 680 -154
rect 700 -163 710 -145
rect 721 -158 736 -154
rect 756 -163 766 -145
rect 797 -134 807 -119
rect 861 -125 871 -119
rect 917 -125 927 -119
rect 812 -163 821 -154
rect 840 -158 855 -154
rect 875 -163 885 -145
rect 896 -158 911 -154
rect 931 -163 941 -145
rect 972 -134 982 -119
rect 1036 -125 1046 -119
rect 1092 -125 1102 -119
rect 987 -163 996 -154
rect 1015 -158 1030 -154
rect 1050 -163 1060 -145
rect 1071 -158 1086 -154
rect 1106 -163 1116 -145
rect 1147 -134 1157 -119
rect 2329 -121 2339 -115
rect 2328 -125 2356 -121
rect 2720 -104 2729 -79
rect 2736 -104 2745 -53
rect 2852 -59 2862 -53
rect 2910 -56 2956 -52
rect 2867 -88 2876 -79
rect 2916 -62 2926 -56
rect 2830 -92 2844 -88
rect 2867 -92 2890 -88
rect 2867 -95 2876 -92
rect 2894 -95 2908 -91
rect 2640 -118 2650 -112
rect 2639 -122 2667 -118
rect 2931 -107 2940 -82
rect 2947 -107 2956 -56
rect 3163 -56 3173 -50
rect 3221 -53 3267 -49
rect 3178 -85 3187 -76
rect 3227 -59 3237 -53
rect 3141 -89 3155 -85
rect 3178 -89 3201 -85
rect 3178 -92 3187 -89
rect 3205 -92 3219 -88
rect 2851 -121 2861 -115
rect 2850 -125 2878 -121
rect 3242 -104 3251 -79
rect 3258 -104 3267 -53
rect 3162 -118 3172 -112
rect 3161 -122 3189 -118
rect 2389 -134 2403 -130
rect 2700 -131 2714 -127
rect 2911 -134 2925 -130
rect 3222 -131 3236 -127
rect 1162 -163 1171 -154
rect 505 -167 614 -163
rect 637 -167 660 -163
rect 680 -167 789 -163
rect 812 -167 835 -163
rect 855 -167 964 -163
rect 987 -167 1010 -163
rect 1030 -167 1139 -163
rect 1162 -167 1185 -163
rect 490 -174 533 -170
rect 490 -305 495 -174
rect 553 -177 563 -167
rect 637 -170 646 -167
rect 693 -174 708 -170
rect 728 -177 738 -167
rect 812 -170 821 -167
rect 537 -203 547 -197
rect 537 -207 563 -203
rect 518 -214 533 -210
rect 553 -217 563 -207
rect 537 -243 547 -237
rect 621 -243 631 -190
rect 868 -174 883 -170
rect 903 -177 913 -167
rect 987 -170 996 -167
rect 712 -203 722 -197
rect 712 -207 738 -203
rect 693 -214 708 -210
rect 728 -217 738 -207
rect 712 -243 722 -237
rect 796 -243 806 -190
rect 1043 -174 1058 -170
rect 1078 -177 1088 -167
rect 1162 -170 1171 -167
rect 887 -203 897 -197
rect 887 -207 913 -203
rect 868 -214 883 -210
rect 903 -217 913 -207
rect 887 -243 897 -237
rect 971 -243 981 -190
rect 1062 -203 1072 -197
rect 1062 -207 1088 -203
rect 1043 -214 1058 -210
rect 1078 -217 1088 -207
rect 1062 -243 1072 -237
rect 1146 -243 1156 -190
rect 2269 -215 2353 -211
rect 2357 -215 2376 -211
rect 2380 -215 2408 -211
rect 2412 -215 2447 -211
rect 2451 -215 2535 -211
rect 2539 -215 2558 -211
rect 2562 -215 2590 -211
rect 2594 -215 2640 -211
rect 2644 -215 2672 -211
rect 2676 -215 2728 -211
rect 2732 -215 2760 -211
rect 2764 -215 2787 -211
rect 2791 -215 2875 -211
rect 2879 -215 2898 -211
rect 2902 -215 2930 -211
rect 2934 -215 2969 -211
rect 2973 -215 3057 -211
rect 3061 -215 3080 -211
rect 3084 -215 3112 -211
rect 3116 -215 3162 -211
rect 3166 -215 3194 -211
rect 3198 -215 3250 -211
rect 3254 -215 3282 -211
rect 2271 -225 2281 -215
rect 2327 -225 2337 -215
rect 509 -247 593 -243
rect 597 -247 616 -243
rect 620 -247 648 -243
rect 652 -247 680 -243
rect 684 -247 768 -243
rect 772 -247 791 -243
rect 795 -247 823 -243
rect 827 -247 855 -243
rect 859 -247 943 -243
rect 947 -247 966 -243
rect 970 -247 998 -243
rect 1002 -247 1030 -243
rect 1034 -247 1118 -243
rect 1122 -247 1141 -243
rect 1145 -247 1173 -243
rect 2250 -258 2265 -254
rect 2285 -263 2295 -245
rect 2306 -258 2321 -254
rect 2341 -263 2351 -245
rect 2382 -234 2392 -215
rect 2453 -225 2463 -215
rect 2509 -225 2519 -215
rect 2397 -263 2406 -254
rect 2432 -258 2447 -254
rect 2467 -263 2477 -245
rect 2488 -258 2503 -254
rect 2523 -263 2533 -245
rect 2564 -234 2574 -215
rect 2646 -221 2656 -215
rect 2626 -254 2640 -250
rect 2579 -263 2588 -254
rect 2660 -257 2670 -241
rect 2640 -261 2676 -257
rect 509 -270 593 -266
rect 597 -270 616 -266
rect 620 -270 648 -266
rect 652 -270 680 -266
rect 684 -270 768 -266
rect 772 -270 791 -266
rect 795 -270 823 -266
rect 827 -270 855 -266
rect 859 -270 943 -266
rect 947 -270 966 -266
rect 970 -270 998 -266
rect 1002 -270 1030 -266
rect 1034 -270 1118 -266
rect 1122 -270 1141 -266
rect 1145 -270 1173 -266
rect 2265 -267 2374 -263
rect 2397 -267 2420 -263
rect 2447 -267 2556 -263
rect 2579 -267 2602 -263
rect 2646 -267 2656 -261
rect 511 -276 521 -270
rect 567 -276 577 -270
rect 490 -309 505 -305
rect 490 -321 495 -309
rect 525 -314 535 -296
rect 546 -309 561 -305
rect 581 -314 591 -296
rect 622 -285 632 -270
rect 686 -276 696 -270
rect 742 -276 752 -270
rect 637 -314 646 -305
rect 665 -309 680 -305
rect 700 -314 710 -296
rect 721 -309 736 -305
rect 756 -314 766 -296
rect 797 -285 807 -270
rect 861 -276 871 -270
rect 917 -276 927 -270
rect 812 -314 821 -305
rect 840 -309 855 -305
rect 875 -314 885 -296
rect 896 -309 911 -305
rect 931 -314 941 -296
rect 972 -285 982 -270
rect 1036 -276 1046 -270
rect 1092 -276 1102 -270
rect 987 -314 996 -305
rect 1015 -309 1030 -305
rect 1050 -314 1060 -296
rect 1071 -309 1086 -305
rect 1106 -314 1116 -296
rect 1147 -285 1157 -270
rect 2278 -274 2293 -270
rect 2313 -277 2323 -267
rect 2397 -270 2406 -267
rect 1162 -314 1171 -305
rect 2460 -274 2475 -270
rect 2495 -277 2505 -267
rect 2579 -270 2588 -267
rect 2297 -303 2307 -297
rect 2297 -307 2323 -303
rect 2278 -314 2293 -310
rect 505 -318 614 -314
rect 637 -318 660 -314
rect 680 -318 789 -314
rect 812 -318 835 -314
rect 855 -318 964 -314
rect 987 -318 1010 -314
rect 1030 -318 1139 -314
rect 1162 -318 1185 -314
rect 2313 -317 2323 -307
rect 490 -325 533 -321
rect 490 -412 495 -325
rect 553 -328 563 -318
rect 637 -321 646 -318
rect 693 -325 708 -321
rect 728 -328 738 -318
rect 812 -321 821 -318
rect 537 -354 547 -348
rect 537 -358 563 -354
rect 518 -365 533 -361
rect 553 -368 563 -358
rect 537 -394 547 -388
rect 621 -394 631 -341
rect 868 -325 883 -321
rect 903 -328 913 -318
rect 987 -321 996 -318
rect 712 -354 722 -348
rect 712 -358 738 -354
rect 693 -365 708 -361
rect 728 -368 738 -358
rect 712 -394 722 -388
rect 796 -394 806 -341
rect 1043 -325 1058 -321
rect 1078 -328 1088 -318
rect 1162 -321 1171 -318
rect 887 -354 897 -348
rect 887 -358 913 -354
rect 868 -365 883 -361
rect 903 -368 913 -358
rect 887 -394 897 -388
rect 971 -394 981 -341
rect 1062 -354 1072 -348
rect 1062 -358 1088 -354
rect 1043 -365 1058 -361
rect 1078 -368 1088 -358
rect 1062 -394 1072 -388
rect 1146 -394 1156 -341
rect 2297 -343 2307 -337
rect 2381 -343 2391 -290
rect 2479 -303 2489 -297
rect 2479 -307 2505 -303
rect 2460 -314 2475 -310
rect 2495 -317 2505 -307
rect 2479 -343 2489 -337
rect 2563 -343 2573 -290
rect 2626 -300 2640 -296
rect 2660 -303 2670 -287
rect 2734 -274 2744 -215
rect 2793 -225 2803 -215
rect 2849 -225 2859 -215
rect 2772 -258 2787 -254
rect 2807 -263 2817 -245
rect 2828 -258 2843 -254
rect 2863 -263 2873 -245
rect 2904 -234 2914 -215
rect 2975 -225 2985 -215
rect 3031 -225 3041 -215
rect 2919 -263 2928 -254
rect 2954 -258 2969 -254
rect 2989 -263 2999 -245
rect 3010 -258 3025 -254
rect 3045 -263 3055 -245
rect 3086 -234 3096 -215
rect 3168 -221 3178 -215
rect 3148 -254 3162 -250
rect 3101 -263 3110 -254
rect 3182 -257 3192 -241
rect 3162 -261 3198 -257
rect 2787 -267 2896 -263
rect 2919 -267 2942 -263
rect 2969 -267 3078 -263
rect 3101 -267 3124 -263
rect 3168 -267 3178 -261
rect 2800 -274 2815 -270
rect 2835 -277 2845 -267
rect 2919 -270 2928 -267
rect 2749 -303 2758 -294
rect 2982 -274 2997 -270
rect 3017 -277 3027 -267
rect 3101 -270 3110 -267
rect 2819 -303 2829 -297
rect 2615 -307 2726 -303
rect 2749 -307 2772 -303
rect 2819 -307 2845 -303
rect 2635 -313 2645 -307
rect 2686 -313 2696 -307
rect 2749 -310 2758 -307
rect 2615 -340 2629 -336
rect 2651 -343 2661 -333
rect 2666 -340 2680 -336
rect 2702 -343 2712 -333
rect 2800 -314 2815 -310
rect 2835 -317 2845 -307
rect 2733 -343 2743 -330
rect 2819 -343 2829 -337
rect 2903 -343 2913 -290
rect 3001 -303 3011 -297
rect 3001 -307 3027 -303
rect 2982 -314 2997 -310
rect 3017 -317 3027 -307
rect 3001 -343 3011 -337
rect 3085 -343 3095 -290
rect 3148 -300 3162 -296
rect 3182 -303 3192 -287
rect 3256 -274 3266 -215
rect 3271 -303 3280 -294
rect 3137 -307 3248 -303
rect 3271 -307 3294 -303
rect 3157 -313 3167 -307
rect 3208 -313 3218 -307
rect 3271 -310 3280 -307
rect 3137 -340 3151 -336
rect 3173 -343 3183 -333
rect 3188 -340 3202 -336
rect 3224 -343 3234 -333
rect 3255 -343 3265 -330
rect 2269 -347 2353 -343
rect 2357 -347 2376 -343
rect 2380 -347 2408 -343
rect 2412 -347 2447 -343
rect 2451 -347 2535 -343
rect 2539 -347 2558 -343
rect 2562 -347 2590 -343
rect 2594 -347 2615 -343
rect 2619 -347 2708 -343
rect 2712 -347 2728 -343
rect 2732 -347 2760 -343
rect 2764 -347 2787 -343
rect 2791 -347 2875 -343
rect 2879 -347 2898 -343
rect 2902 -347 2930 -343
rect 2934 -347 2969 -343
rect 2973 -347 3057 -343
rect 3061 -347 3080 -343
rect 3084 -347 3112 -343
rect 3116 -347 3137 -343
rect 3141 -347 3230 -343
rect 3234 -347 3250 -343
rect 3254 -347 3282 -343
rect 2328 -357 2356 -353
rect 2387 -357 2434 -353
rect 2639 -354 2667 -350
rect 2698 -354 2745 -350
rect 2330 -363 2340 -357
rect 2393 -363 2403 -357
rect 2345 -392 2354 -383
rect 509 -398 593 -394
rect 597 -398 616 -394
rect 620 -398 648 -394
rect 652 -398 680 -394
rect 684 -398 768 -394
rect 772 -398 791 -394
rect 795 -398 823 -394
rect 827 -398 855 -394
rect 859 -398 943 -394
rect 947 -398 966 -394
rect 970 -398 998 -394
rect 1002 -398 1030 -394
rect 1034 -398 1118 -394
rect 1122 -398 1141 -394
rect 1145 -398 1173 -394
rect 1177 -398 1197 -394
rect 2308 -396 2322 -392
rect 2345 -396 2368 -392
rect 2372 -396 2385 -392
rect 2345 -399 2354 -396
rect 490 -417 1020 -412
rect 2408 -408 2417 -383
rect 2424 -408 2434 -357
rect 2641 -360 2651 -354
rect 2704 -360 2714 -354
rect 2656 -389 2665 -380
rect 2619 -393 2633 -389
rect 2656 -393 2679 -389
rect 2683 -393 2696 -389
rect 2656 -396 2665 -393
rect 2329 -425 2339 -419
rect 2328 -429 2356 -425
rect 2719 -405 2728 -380
rect 2735 -405 2745 -354
rect 2850 -357 2878 -353
rect 2909 -357 2956 -353
rect 3161 -354 3189 -350
rect 3220 -354 3267 -350
rect 2852 -363 2862 -357
rect 2915 -363 2925 -357
rect 2867 -392 2876 -383
rect 2830 -396 2844 -392
rect 2867 -396 2890 -392
rect 2894 -396 2907 -392
rect 2867 -399 2876 -396
rect 2640 -422 2650 -416
rect 2639 -426 2667 -422
rect 2930 -408 2939 -383
rect 2946 -408 2956 -357
rect 3163 -360 3173 -354
rect 3226 -360 3236 -354
rect 3178 -389 3187 -380
rect 3141 -393 3155 -389
rect 3178 -393 3201 -389
rect 3205 -393 3218 -389
rect 3178 -396 3187 -393
rect 2851 -425 2861 -419
rect 2388 -435 2402 -431
rect 2699 -432 2713 -428
rect 2850 -429 2878 -425
rect 3241 -405 3250 -380
rect 3257 -405 3267 -354
rect 3162 -422 3172 -416
rect 3161 -426 3189 -422
rect 2328 -439 2356 -435
rect 2639 -436 2667 -432
rect 2910 -435 2924 -431
rect 3221 -432 3235 -428
rect 632 -445 660 -441
rect 691 -445 738 -441
rect 773 -445 801 -441
rect 832 -445 879 -441
rect 917 -445 1112 -441
rect 1116 -445 1134 -441
rect 1138 -445 1166 -441
rect 2330 -445 2340 -439
rect 2388 -442 2434 -438
rect 634 -451 644 -445
rect 697 -451 707 -445
rect 649 -480 658 -471
rect 612 -484 626 -480
rect 649 -484 672 -480
rect 675 -484 689 -480
rect 649 -487 658 -484
rect 712 -496 721 -471
rect 728 -496 738 -445
rect 775 -451 785 -445
rect 838 -451 848 -445
rect 790 -480 799 -471
rect 753 -484 767 -480
rect 790 -484 813 -480
rect 816 -484 830 -480
rect 790 -487 799 -484
rect 633 -513 643 -507
rect 632 -517 660 -513
rect 853 -496 862 -471
rect 869 -496 879 -445
rect 919 -451 929 -445
rect 975 -451 985 -445
rect 1031 -451 1041 -445
rect 1087 -451 1097 -445
rect 898 -484 913 -480
rect 933 -489 943 -471
rect 954 -484 969 -480
rect 989 -489 999 -471
rect 1010 -484 1025 -480
rect 1045 -489 1055 -471
rect 1066 -484 1081 -480
rect 1101 -489 1111 -471
rect 1139 -460 1149 -445
rect 2345 -474 2354 -465
rect 2394 -448 2404 -442
rect 2308 -478 2322 -474
rect 2345 -478 2368 -474
rect 1154 -489 1163 -480
rect 2345 -481 2354 -478
rect 2372 -481 2386 -477
rect 913 -493 1131 -489
rect 1154 -493 1177 -489
rect 774 -513 784 -507
rect 773 -517 801 -513
rect 926 -500 941 -496
rect 961 -503 971 -493
rect 1154 -496 1163 -493
rect 692 -523 706 -519
rect 833 -523 847 -519
rect 2409 -493 2418 -468
rect 2425 -493 2434 -442
rect 2641 -442 2651 -436
rect 2699 -439 2745 -435
rect 2850 -439 2878 -435
rect 3161 -436 3189 -432
rect 2656 -471 2665 -462
rect 2705 -445 2715 -439
rect 2619 -475 2633 -471
rect 2656 -475 2679 -471
rect 2656 -478 2665 -475
rect 2683 -478 2697 -474
rect 1234 -510 1485 -506
rect 2329 -507 2339 -501
rect 1236 -516 1246 -510
rect 1292 -516 1302 -510
rect 1348 -516 1358 -510
rect 1404 -516 1414 -510
rect 1459 -516 1469 -510
rect 2328 -511 2356 -507
rect 2720 -490 2729 -465
rect 2736 -490 2745 -439
rect 2852 -445 2862 -439
rect 2910 -442 2956 -438
rect 2867 -474 2876 -465
rect 2916 -448 2926 -442
rect 2830 -478 2844 -474
rect 2867 -478 2890 -474
rect 2867 -481 2876 -478
rect 2894 -481 2908 -477
rect 2640 -504 2650 -498
rect 2639 -508 2667 -504
rect 2931 -493 2940 -468
rect 2947 -493 2956 -442
rect 3163 -442 3173 -436
rect 3221 -439 3267 -435
rect 3178 -471 3187 -462
rect 3227 -445 3237 -439
rect 3141 -475 3155 -471
rect 3178 -475 3201 -471
rect 3178 -478 3187 -475
rect 3205 -478 3219 -474
rect 2851 -507 2861 -501
rect 2850 -511 2878 -507
rect 3242 -490 3251 -465
rect 3258 -490 3267 -439
rect 3162 -504 3172 -498
rect 3161 -508 3189 -504
rect 632 -527 660 -523
rect 634 -533 644 -527
rect 692 -530 738 -526
rect 773 -527 801 -523
rect 649 -562 658 -553
rect 698 -536 708 -530
rect 612 -566 626 -562
rect 649 -566 672 -562
rect 649 -569 658 -566
rect 676 -569 690 -565
rect 713 -581 722 -556
rect 729 -581 738 -530
rect 775 -533 785 -527
rect 833 -530 879 -526
rect 790 -562 799 -553
rect 839 -536 849 -530
rect 753 -566 767 -562
rect 790 -566 813 -562
rect 790 -569 799 -566
rect 817 -569 831 -565
rect 633 -595 643 -589
rect 632 -599 660 -595
rect 854 -581 863 -556
rect 870 -581 879 -530
rect 945 -529 955 -523
rect 945 -533 971 -529
rect 926 -540 941 -536
rect 961 -543 971 -533
rect 945 -569 955 -563
rect 945 -573 971 -569
rect 926 -580 941 -576
rect 774 -595 784 -589
rect 773 -599 801 -595
rect 961 -583 971 -573
rect 693 -608 707 -604
rect 834 -608 848 -604
rect 945 -608 955 -603
rect 945 -612 971 -608
rect 926 -619 941 -615
rect 961 -622 971 -612
rect 632 -626 660 -622
rect 691 -626 738 -622
rect 773 -626 801 -622
rect 832 -626 879 -622
rect 634 -632 644 -626
rect 697 -632 707 -626
rect 649 -661 658 -652
rect 612 -665 626 -661
rect 649 -665 672 -661
rect 675 -665 689 -661
rect 649 -668 658 -665
rect 712 -677 721 -652
rect 728 -677 738 -626
rect 775 -632 785 -626
rect 838 -632 848 -626
rect 790 -661 799 -652
rect 753 -665 767 -661
rect 790 -665 813 -661
rect 816 -665 830 -661
rect 790 -668 799 -665
rect 633 -694 643 -688
rect 632 -698 660 -694
rect 853 -677 862 -652
rect 869 -677 879 -626
rect 945 -647 955 -642
rect 1138 -647 1148 -516
rect 2389 -520 2403 -516
rect 2700 -517 2714 -513
rect 2911 -520 2925 -516
rect 3222 -517 3236 -513
rect 1215 -549 1230 -545
rect 1250 -554 1260 -536
rect 1271 -549 1286 -545
rect 1306 -554 1316 -536
rect 1327 -549 1342 -545
rect 1362 -554 1372 -536
rect 1383 -549 1398 -545
rect 1418 -554 1428 -536
rect 1438 -549 1453 -545
rect 1473 -554 1483 -536
rect 1230 -558 1489 -554
rect 1243 -565 1258 -561
rect 1278 -568 1288 -558
rect 1596 -581 1680 -577
rect 1684 -581 1703 -577
rect 1707 -581 1735 -577
rect 1739 -581 1762 -577
rect 1766 -581 1850 -577
rect 1854 -581 1873 -577
rect 1877 -581 1905 -577
rect 1909 -581 1932 -577
rect 1936 -581 2020 -577
rect 2024 -581 2043 -577
rect 2047 -581 2075 -577
rect 2079 -581 2102 -577
rect 2106 -581 2190 -577
rect 2194 -581 2213 -577
rect 2217 -581 2245 -577
rect 1598 -587 1608 -581
rect 1654 -587 1664 -581
rect 1262 -594 1272 -588
rect 1262 -598 1288 -594
rect 1243 -605 1258 -601
rect 1278 -608 1288 -598
rect 1577 -620 1592 -616
rect 1612 -625 1622 -607
rect 1633 -620 1648 -616
rect 1668 -625 1678 -607
rect 1709 -596 1719 -581
rect 1768 -587 1778 -581
rect 1824 -587 1834 -581
rect 1724 -625 1733 -616
rect 1747 -620 1762 -616
rect 1782 -625 1792 -607
rect 1803 -620 1818 -616
rect 1838 -625 1848 -607
rect 1879 -596 1889 -581
rect 1938 -587 1948 -581
rect 1994 -587 2004 -581
rect 1894 -625 1903 -616
rect 1917 -620 1932 -616
rect 1952 -625 1962 -607
rect 1973 -620 1988 -616
rect 2008 -625 2018 -607
rect 2049 -596 2059 -581
rect 2108 -587 2118 -581
rect 2164 -587 2174 -581
rect 2064 -625 2073 -616
rect 2087 -620 2102 -616
rect 2122 -625 2132 -607
rect 2143 -620 2158 -616
rect 2178 -625 2188 -607
rect 2219 -596 2229 -581
rect 2234 -625 2243 -616
rect 1262 -634 1272 -628
rect 1592 -629 1701 -625
rect 1724 -629 1747 -625
rect 1762 -629 1871 -625
rect 1894 -629 1917 -625
rect 1932 -629 2041 -625
rect 2064 -629 2087 -625
rect 2102 -629 2211 -625
rect 2234 -629 2257 -625
rect 1262 -638 1288 -634
rect 1605 -636 1620 -632
rect 1243 -645 1258 -641
rect 917 -651 1113 -647
rect 1117 -651 1134 -647
rect 1138 -651 1166 -647
rect 1278 -648 1288 -638
rect 1640 -639 1650 -629
rect 1724 -632 1733 -629
rect 947 -662 1031 -658
rect 1072 -662 1097 -658
rect 1101 -662 1129 -658
rect 1133 -662 1169 -658
rect 774 -694 784 -688
rect 773 -698 801 -694
rect 949 -668 959 -662
rect 1005 -668 1015 -662
rect 1103 -668 1113 -662
rect 1775 -636 1790 -632
rect 1810 -639 1820 -629
rect 1894 -632 1903 -629
rect 1624 -665 1634 -659
rect 1262 -673 1272 -668
rect 1624 -669 1650 -665
rect 1262 -677 1288 -673
rect 1605 -676 1620 -672
rect 1243 -684 1258 -680
rect 1278 -687 1288 -677
rect 1640 -679 1650 -669
rect 692 -704 706 -700
rect 833 -704 847 -700
rect 928 -701 943 -697
rect 632 -708 660 -704
rect 634 -714 644 -708
rect 692 -711 738 -707
rect 773 -708 801 -704
rect 963 -706 973 -688
rect 984 -701 999 -697
rect 1019 -706 1029 -688
rect 1083 -701 1097 -697
rect 1117 -704 1127 -688
rect 649 -743 658 -734
rect 698 -717 708 -711
rect 612 -747 626 -743
rect 649 -747 672 -743
rect 649 -750 658 -747
rect 676 -750 690 -746
rect 713 -762 722 -737
rect 729 -762 738 -711
rect 775 -714 785 -708
rect 833 -711 879 -707
rect 943 -710 1035 -706
rect 1097 -708 1133 -704
rect 1624 -705 1634 -699
rect 1708 -705 1718 -652
rect 1945 -636 1960 -632
rect 1980 -639 1990 -629
rect 2064 -632 2073 -629
rect 1794 -665 1804 -659
rect 1794 -669 1820 -665
rect 1775 -676 1790 -672
rect 1810 -679 1820 -669
rect 1794 -705 1804 -699
rect 1878 -705 1888 -652
rect 2115 -636 2130 -632
rect 2150 -639 2160 -629
rect 2234 -632 2243 -629
rect 1964 -665 1974 -659
rect 1964 -669 1990 -665
rect 1945 -676 1960 -672
rect 1980 -679 1990 -669
rect 1964 -705 1974 -699
rect 2048 -705 2058 -652
rect 2134 -665 2144 -659
rect 2134 -669 2160 -665
rect 2115 -676 2130 -672
rect 2150 -679 2160 -669
rect 2134 -705 2144 -699
rect 2218 -705 2228 -652
rect 790 -743 799 -734
rect 839 -717 849 -711
rect 753 -747 767 -743
rect 790 -747 813 -743
rect 790 -750 799 -747
rect 817 -750 831 -746
rect 633 -776 643 -770
rect 632 -780 660 -776
rect 854 -762 863 -737
rect 870 -762 879 -711
rect 956 -717 971 -713
rect 991 -720 1001 -710
rect 1103 -714 1113 -708
rect 1262 -712 1272 -707
rect 1596 -709 1680 -705
rect 1684 -709 1703 -705
rect 1707 -709 1735 -705
rect 1739 -709 1762 -705
rect 1766 -709 1850 -705
rect 1854 -709 1873 -705
rect 1877 -709 1905 -705
rect 1909 -709 1932 -705
rect 1936 -709 2020 -705
rect 2024 -709 2043 -705
rect 2047 -709 2075 -705
rect 2079 -709 2102 -705
rect 2106 -709 2190 -705
rect 2194 -709 2213 -705
rect 2217 -709 2245 -705
rect 1262 -716 1288 -712
rect 1243 -723 1258 -719
rect 1278 -726 1288 -716
rect 975 -746 985 -740
rect 975 -750 1001 -746
rect 1083 -747 1097 -743
rect 1117 -750 1127 -734
rect 956 -757 971 -753
rect 991 -760 1001 -750
rect 1072 -754 1169 -750
rect 1262 -751 1272 -746
rect 774 -776 784 -770
rect 773 -780 801 -776
rect 1092 -760 1102 -754
rect 1143 -760 1153 -754
rect 1234 -755 1485 -751
rect 693 -789 707 -785
rect 834 -789 848 -785
rect 975 -786 985 -780
rect 947 -790 1031 -786
rect 1072 -787 1086 -783
rect 1108 -790 1118 -780
rect 1123 -787 1137 -783
rect 1159 -790 1169 -780
rect 1076 -794 1165 -790
rect 632 -807 772 -803
rect 840 -806 1036 -802
rect 1132 -806 1328 -802
rect 634 -813 644 -807
rect 690 -813 700 -807
rect 746 -813 756 -807
rect 842 -812 852 -806
rect 898 -812 908 -806
rect 954 -812 964 -806
rect 1010 -812 1020 -806
rect 1134 -812 1144 -806
rect 1190 -812 1200 -806
rect 1246 -812 1256 -806
rect 1302 -812 1312 -806
rect 613 -846 628 -842
rect 648 -851 658 -833
rect 669 -846 684 -842
rect 704 -851 714 -833
rect 725 -846 740 -842
rect 760 -851 770 -833
rect 821 -845 836 -841
rect 856 -850 866 -832
rect 877 -845 892 -841
rect 912 -850 922 -832
rect 933 -845 948 -841
rect 968 -850 978 -832
rect 989 -845 1004 -841
rect 1024 -850 1034 -832
rect 1113 -845 1128 -841
rect 1148 -850 1158 -832
rect 1169 -845 1184 -841
rect 1204 -850 1214 -832
rect 1225 -845 1240 -841
rect 1260 -850 1270 -832
rect 1281 -845 1296 -841
rect 1316 -850 1326 -832
rect 628 -855 776 -851
rect 836 -854 1040 -850
rect 1128 -854 1332 -850
rect 641 -862 656 -858
rect 676 -865 686 -855
rect 849 -861 864 -857
rect 884 -864 894 -854
rect 1141 -861 1156 -857
rect 1176 -864 1186 -854
rect 1414 -884 1498 -880
rect 1502 -884 1521 -880
rect 1525 -884 1553 -880
rect 660 -891 670 -885
rect 868 -890 878 -884
rect 1160 -890 1170 -884
rect 1416 -890 1426 -884
rect 1472 -890 1482 -884
rect 660 -895 686 -891
rect 868 -894 894 -890
rect 1160 -894 1186 -890
rect 641 -902 656 -898
rect 676 -905 686 -895
rect 849 -901 864 -897
rect 884 -904 894 -894
rect 1141 -901 1156 -897
rect 1176 -904 1186 -894
rect 1395 -923 1410 -919
rect 660 -931 670 -925
rect 868 -930 878 -924
rect 1160 -930 1170 -924
rect 1430 -928 1440 -910
rect 1451 -923 1466 -919
rect 1486 -928 1496 -910
rect 1527 -899 1537 -884
rect 1542 -928 1551 -919
rect 660 -935 686 -931
rect 868 -934 894 -930
rect 1160 -934 1186 -930
rect 1410 -932 1519 -928
rect 1542 -932 1565 -928
rect 641 -942 656 -938
rect 676 -945 686 -935
rect 849 -941 864 -937
rect 884 -944 894 -934
rect 1141 -941 1156 -937
rect 1176 -944 1186 -934
rect 1423 -939 1438 -935
rect 1458 -942 1468 -932
rect 1542 -935 1551 -932
rect 660 -970 670 -965
rect 868 -969 878 -964
rect 1160 -969 1170 -964
rect 1442 -968 1452 -962
rect 632 -974 772 -970
rect 868 -973 894 -969
rect 1160 -973 1186 -969
rect 1442 -972 1468 -968
rect 849 -980 864 -976
rect 884 -983 894 -973
rect 1141 -980 1156 -976
rect 1176 -983 1186 -973
rect 1423 -979 1438 -975
rect 1458 -982 1468 -972
rect 868 -1008 878 -1003
rect 1160 -1008 1170 -1003
rect 1442 -1008 1452 -1002
rect 1526 -1008 1536 -955
rect 840 -1012 1036 -1008
rect 1132 -1012 1328 -1008
rect 1414 -1012 1498 -1008
rect 1502 -1012 1521 -1008
rect 1525 -1012 1553 -1008
<< metal2 >>
rect 622 555 627 597
rect 797 555 802 597
rect 972 555 977 597
rect 622 296 627 383
rect 797 296 802 383
rect 972 296 977 383
rect 766 222 771 291
rect 1320 244 1325 304
rect 1495 244 1500 304
rect 1670 244 1675 304
rect 942 79 985 83
rect 981 50 985 79
rect 969 46 992 50
rect 969 -6 973 46
rect 1033 -6 1037 6
rect 969 -10 1037 -6
rect 1320 -23 1325 72
rect 1495 -23 1500 72
rect 1670 -23 1675 72
<< m123contact >>
rect 622 597 627 602
rect 622 550 627 555
rect 797 597 802 602
rect 797 550 802 555
rect 972 597 977 602
rect 972 550 977 555
rect 622 383 627 388
rect 797 383 802 388
rect 622 291 627 296
rect 766 291 771 296
rect 797 291 802 296
rect 972 383 977 388
rect 972 291 977 296
rect 1320 304 1325 309
rect 1320 239 1325 244
rect 1495 304 1500 309
rect 1495 239 1500 244
rect 1670 304 1675 309
rect 1670 239 1675 244
rect 766 217 771 222
rect 992 92 997 97
rect 767 79 772 84
rect 937 79 942 84
rect 1320 72 1325 77
rect 992 46 997 51
rect 981 6 986 11
rect 1033 6 1038 11
rect 1320 -28 1325 -23
rect 1495 72 1500 77
rect 1495 -28 1500 -23
rect 1670 72 1675 77
rect 1670 -28 1675 -23
<< metal3 >>
rect 977 92 992 96
rect 772 79 780 83
rect 776 -12 780 79
rect 977 10 981 92
rect 973 6 981 10
rect 973 -12 977 6
rect 776 -16 977 -12
<< labels >>
rlabel metal1 558 -1 965 3 1 Gnd
rlabel metal1 526 265 933 269 5 VDD
rlabel metal1 542 170 560 174 1 S1
rlabel metal1 584 170 602 174 1 S1not
rlabel metal1 543 32 560 36 1 S0
rlabel metal1 585 32 602 36 1 S0not
rlabel metal1 601 226 620 230 1 S1
rlabel metal1 629 210 648 214 1 S1
rlabel metal1 657 226 676 230 1 S0
rlabel metal1 629 170 648 174 1 S0
rlabel metal1 752 217 771 221 1 D3
rlabel metal1 771 226 790 230 1 S1
rlabel metal1 799 210 818 214 1 S1
rlabel metal1 827 226 846 230 1 S0not
rlabel metal1 799 170 818 174 1 S0not
rlabel metal1 922 217 941 221 1 D2
rlabel metal1 601 88 620 92 1 S1not
rlabel metal1 629 72 648 76 1 S1not
rlabel metal1 657 88 676 92 1 S0
rlabel metal1 629 32 648 36 1 S0
rlabel metal1 752 79 771 83 1 D1
rlabel metal1 771 88 790 92 1 S1not
rlabel metal1 799 72 818 76 1 S1not
rlabel metal1 827 88 846 92 1 S0not
rlabel metal1 799 32 818 36 1 S0not
rlabel metal1 922 79 941 83 1 D0
rlabel metal1 982 131 1131 135 5 VDD
rlabel metal1 982 -1 1131 3 1 Gnd
rlabel metal1 993 92 1011 96 1 D1
rlabel metal1 982 6 1000 10 1 D1
rlabel metal1 1121 39 1139 43 1 DAS
rlabel metal1 518 -365 537 -361 1 B3
rlabel metal1 693 -365 712 -361 1 B2
rlabel metal1 868 -365 887 -361 1 B1
rlabel metal1 1043 -365 1062 -361 1 B0
rlabel metal1 1071 -309 1090 -305 1 B0
rlabel metal1 896 -309 915 -305 1 B1
rlabel metal1 721 -309 740 -305 1 B2
rlabel metal1 546 -309 565 -305 1 B3
rlabel metal1 505 -398 1197 -394 1 Gnd
rlabel metal1 505 -247 1177 -243 1 Gnd
rlabel metal1 505 -270 1177 -266 1 VDD
rlabel metal1 505 -119 1177 -115 5 VDD
rlabel metal1 518 -214 537 -210 1 A3
rlabel metal1 693 -214 712 -210 1 A2
rlabel metal1 868 -214 887 -210 1 A1
rlabel metal1 1043 -214 1062 -210 1 A0
rlabel metal1 1071 -158 1090 -154 1 A0
rlabel metal1 896 -158 915 -154 1 A1
rlabel metal1 721 -158 740 -154 1 A2
rlabel metal1 546 -158 565 -154 1 A3
rlabel metal1 490 -158 509 -154 1 D2
rlabel metal1 518 -174 537 -170 1 D2
rlabel metal1 665 -158 684 -154 1 D2
rlabel metal1 693 -174 712 -170 1 D2
rlabel metal1 840 -158 859 -154 1 D2
rlabel metal1 868 -174 887 -170 1 D2
rlabel metal1 1015 -158 1034 -154 1 D2
rlabel metal1 1043 -174 1062 -170 1 D2
rlabel metal1 641 -167 660 -163 1 COA3
rlabel metal1 816 -167 835 -163 1 COA2
rlabel metal1 991 -167 1010 -163 1 COA1
rlabel metal1 1166 -167 1185 -163 1 COA0
rlabel metal1 1166 -318 1185 -314 1 COB0
rlabel metal1 991 -318 1010 -314 1 COB1
rlabel metal1 816 -318 835 -314 1 COB2
rlabel metal1 641 -318 660 -314 1 COB3
rlabel metal1 490 -309 509 -305 1 D2
rlabel metal1 518 -325 537 -321 1 D2
rlabel metal1 665 -309 684 -305 1 D2
rlabel metal1 693 -325 712 -321 1 D2
rlabel metal1 840 -309 859 -305 1 D2
rlabel metal1 868 -325 887 -321 1 D2
rlabel metal1 1015 -309 1034 -305 1 D2
rlabel metal1 1043 -325 1062 -321 1 D2
rlabel metal1 2265 39 2764 43 1 Gnd
rlabel metal1 2324 -43 2360 -39 1 Gnd
rlabel metal1 2324 -53 2360 -49 1 VDD
rlabel metal1 2324 -125 2360 -121 1 Gnd
rlabel metal1 2324 29 2360 33 1 VDD
rlabel metal1 2635 32 2671 36 1 VDD
rlabel metal1 2635 -50 2671 -46 1 VDD
rlabel metal1 2635 -40 2671 -36 1 Gnd
rlabel metal1 2635 -122 2671 -118 1 Gnd
rlabel metal1 2787 39 3286 43 1 Gnd
rlabel metal1 2846 -43 2882 -39 1 Gnd
rlabel metal1 2846 -53 2882 -49 1 VDD
rlabel metal1 2846 -125 2882 -121 1 Gnd
rlabel metal1 2846 29 2882 33 1 VDD
rlabel metal1 3157 32 3193 36 1 VDD
rlabel metal1 3157 -50 3193 -46 1 VDD
rlabel metal1 3157 -40 3193 -36 1 Gnd
rlabel metal1 3157 -122 3193 -118 1 Gnd
rlabel metal1 2754 -307 2772 -303 1 C
rlabel metal1 2265 -347 2764 -343 1 Gnd
rlabel metal1 2324 -429 2360 -425 1 Gnd
rlabel metal1 2324 -439 2360 -435 1 VDD
rlabel metal1 2324 -511 2360 -507 1 Gnd
rlabel metal1 2324 -357 2360 -353 1 VDD
rlabel metal1 2635 -354 2671 -350 1 VDD
rlabel metal1 2635 -436 2671 -432 1 VDD
rlabel metal1 2635 -426 2671 -422 1 Gnd
rlabel metal1 2635 -508 2671 -504 1 Gnd
rlabel metal1 2787 -347 3286 -343 1 Gnd
rlabel metal1 2846 -429 2882 -425 1 Gnd
rlabel metal1 2846 -439 2882 -435 1 VDD
rlabel metal1 2846 -511 2882 -507 1 Gnd
rlabel metal1 2846 -357 2882 -353 1 VDD
rlabel metal1 3157 -354 3193 -350 1 VDD
rlabel metal1 3157 -436 3193 -432 1 VDD
rlabel metal1 3157 -426 3193 -422 1 Gnd
rlabel metal1 3157 -508 3193 -504 1 Gnd
rlabel metal1 2265 171 2615 175 1 VDD
rlabel metal1 2787 171 3137 175 1 VDD
rlabel metal1 2265 -215 2615 -211 1 VDD
rlabel metal1 2787 -215 3137 -211 1 VDD
rlabel metal1 2250 -258 2269 -254 1 ASA3
rlabel metal1 2278 -274 2297 -270 1 ASA3
rlabel metal1 2306 -258 2325 -254 1 xorB3
rlabel metal1 2278 -314 2297 -310 1 xorB3
rlabel metal1 2401 -267 2420 -263 1 FA3C2
rlabel metal1 2432 -258 2451 -254 1 FA3S1
rlabel metal1 2488 -258 2507 -254 1 C2
rlabel metal1 2460 -274 2479 -270 1 FA3S1
rlabel metal1 2460 -314 2479 -310 1 C2
rlabel metal1 2583 -267 2602 -263 1 FA3C1
rlabel metal1 2308 -396 2326 -392 1 ASA3
rlabel metal1 2350 -396 2368 -392 1 ASA3not
rlabel metal1 2372 -396 2389 -392 1 xorB3
rlabel metal1 2308 -478 2326 -474 1 xorB3
rlabel metal1 2350 -478 2368 -474 1 xorB3not
rlabel metal1 2388 -435 2406 -431 1 xorB3not
rlabel metal1 2372 -481 2390 -477 1 xorB3not
rlabel metal1 2389 -520 2407 -516 1 xorB3
rlabel metal1 2408 -408 2417 -389 1 ASA3
rlabel metal1 2409 -493 2418 -474 1 ASA3not
rlabel metal1 2424 -408 2434 -353 1 FA3S1
rlabel metal1 2425 -493 2434 -438 1 FA3S1
rlabel metal1 2619 -393 2637 -389 1 FA3S1
rlabel metal1 2661 -393 2679 -389 1 FA3S1not
rlabel metal1 2619 -475 2637 -471 1 C2
rlabel metal1 2661 -475 2679 -471 1 C2not
rlabel metal1 2719 -405 2728 -386 1 C2
rlabel metal1 2720 -490 2729 -471 1 C2not
rlabel metal1 2735 -405 2745 -350 1 OUT_AS3
rlabel metal1 2736 -490 2745 -435 1 OUT_AS3
rlabel metal1 2683 -393 2700 -389 1 FA3S1
rlabel metal1 2699 -432 2717 -428 1 FA3S1not
rlabel metal1 2683 -478 2701 -474 1 FA3S1not
rlabel metal1 2700 -517 2718 -513 1 FA3S1
rlabel metal1 2626 -254 2644 -250 1 FA3C1
rlabel metal1 2626 -300 2644 -296 1 FA3C2
rlabel metal1 2615 -340 2633 -336 1 FA3C1
rlabel metal1 2666 -340 2684 -336 1 FA3C2
rlabel metal1 2772 -258 2791 -254 1 ASA2
rlabel metal1 2800 -274 2819 -270 1 ASA2
rlabel metal1 2830 -396 2848 -392 1 ASA2
rlabel metal1 2872 -396 2890 -392 1 ASA2not
rlabel metal1 2828 -258 2847 -254 1 xorB2
rlabel metal1 2800 -314 2819 -310 1 xorB2
rlabel metal1 2830 -478 2848 -474 1 xorB2
rlabel metal1 2872 -478 2890 -474 1 xorB2not
rlabel metal1 2910 -435 2928 -431 1 xorB2not
rlabel metal1 2894 -481 2912 -477 1 xorB2not
rlabel metal1 2894 -396 2911 -392 1 xorB2
rlabel metal1 2911 -520 2929 -516 1 xorB2
rlabel metal1 2930 -408 2939 -389 1 ASA2
rlabel metal1 2931 -493 2940 -474 1 ASA2not
rlabel metal1 2947 -493 2956 -438 1 FA2S1
rlabel metal1 2946 -408 2956 -353 1 FA2S1
rlabel metal1 3141 -393 3159 -389 1 FA2S1
rlabel metal1 3183 -393 3201 -389 1 FA2S1not
rlabel metal1 3141 -475 3159 -471 1 C1
rlabel metal1 3183 -475 3201 -471 1 C1not
rlabel metal1 3241 -405 3250 -386 1 C1
rlabel metal1 3242 -490 3251 -471 1 C1not
rlabel metal1 3205 -393 3222 -389 1 FA2S1
rlabel metal1 3205 -478 3223 -474 1 FA2S1not
rlabel metal1 3221 -432 3239 -428 1 FA2S1not
rlabel metal1 3222 -517 3240 -513 1 FA2S1
rlabel metal1 3258 -490 3267 -435 1 OUT_AS2
rlabel metal1 3257 -405 3267 -350 1 OUT_AS2
rlabel metal1 2923 -267 2942 -263 1 FA2C2
rlabel metal1 2954 -258 2973 -254 1 FA2S1
rlabel metal1 2982 -274 3001 -270 1 FA2S1
rlabel metal1 3105 -267 3124 -263 1 FA2C1
rlabel metal1 3148 -254 3166 -250 1 FA2C1
rlabel metal1 3137 -340 3155 -336 1 FA2C1
rlabel metal1 3148 -300 3166 -296 1 FA2C2
rlabel metal1 3188 -340 3206 -336 1 FA2C2
rlabel metal1 3010 -258 3029 -254 1 C1
rlabel metal1 2982 -314 3001 -310 1 C1
rlabel metal1 3276 -307 3294 -303 1 C2
rlabel metal1 2772 128 2791 132 1 ASA1
rlabel metal1 2800 112 2819 116 1 ASA1
rlabel metal1 2830 -10 2848 -6 1 ASA1
rlabel metal1 2872 -10 2890 -6 1 ASA1not
rlabel metal1 2930 -22 2939 -3 1 ASA1
rlabel metal1 2931 -107 2940 -88 1 ASA1not
rlabel metal1 2946 -22 2956 33 1 FA1S1
rlabel metal1 2947 -107 2956 -52 1 FA1S1
rlabel metal1 2828 128 2847 132 1 xorB1
rlabel metal1 2800 72 2819 76 1 xorB1
rlabel metal1 2830 -92 2848 -88 1 xorB1
rlabel metal1 2894 -10 2911 -6 1 xorB1
rlabel metal1 2911 -134 2929 -130 1 xorB1
rlabel metal1 2872 -92 2890 -88 1 xorB1not
rlabel metal1 2910 -49 2928 -45 1 xorB1not
rlabel metal1 2894 -95 2912 -91 1 xorB1not
rlabel metal1 2923 119 2942 123 1 FA1C2
rlabel metal1 2954 128 2973 132 1 FA1S1
rlabel metal1 2982 112 3001 116 1 FA1S1
rlabel metal1 3010 128 3029 132 1 C0
rlabel metal1 2982 72 3001 76 1 C0
rlabel metal1 3105 119 3124 123 1 FA1C1
rlabel metal1 3141 -7 3159 -3 1 FA1S1
rlabel metal1 3222 -131 3240 -127 1 FA1S1
rlabel metal1 3183 -7 3201 -3 1 FA1S1not
rlabel metal1 3141 -89 3159 -85 1 C0
rlabel metal1 3183 -89 3201 -85 1 C0not
rlabel metal1 3205 -7 3222 -3 1 FA1S1
rlabel metal1 3221 -46 3239 -42 1 FA1S1not
rlabel metal1 3205 -92 3223 -88 1 FA1S1not
rlabel metal1 3241 -19 3250 0 1 C0
rlabel metal1 3242 -104 3251 -85 1 C0not
rlabel metal1 3258 -104 3267 -49 1 OUT_AS1
rlabel metal1 3257 -19 3267 36 1 OUT_AS1
rlabel metal1 3148 132 3166 136 1 FA1C1
rlabel metal1 3148 86 3166 90 1 FA1C2
rlabel metal1 3188 46 3206 50 1 FA1C2
rlabel metal1 3137 46 3155 50 1 FA1C1
rlabel metal1 3276 79 3294 83 1 C1
rlabel metal1 2250 128 2269 132 1 ASA0
rlabel metal1 2278 112 2297 116 1 ASA0
rlabel metal1 2308 -10 2326 -6 1 ASA0
rlabel metal1 2350 -10 2368 -6 1 ASA0not
rlabel metal1 2278 72 2297 76 1 xorB0
rlabel metal1 2306 128 2325 132 1 xorB0
rlabel metal1 2308 -92 2326 -88 1 xorB0
rlabel metal1 2350 -92 2368 -88 1 xorB0not
rlabel metal1 2372 -95 2390 -91 1 xorB0not
rlabel metal1 2388 -49 2406 -45 1 xorB0not
rlabel metal1 2372 -10 2389 -6 1 xorB0
rlabel metal1 2389 -134 2407 -130 1 xorB0
rlabel metal1 2408 -22 2417 -3 1 ASA0
rlabel metal1 2409 -107 2418 -88 1 ASA0not
rlabel metal1 2425 -107 2434 -52 1 FA0S1
rlabel metal1 2424 -22 2434 33 1 FA0S1
rlabel metal1 2401 119 2420 123 1 FA0C2
rlabel metal1 2432 128 2451 132 1 FA0S1
rlabel metal1 2460 112 2479 116 1 FA0S1
rlabel metal1 2488 128 2507 132 1 D1
rlabel metal1 2460 72 2479 76 1 D1
rlabel metal1 2583 119 2602 123 1 FA0C1
rlabel metal1 2626 132 2644 136 1 FA0C1
rlabel metal1 2615 46 2633 50 1 FA0C1
rlabel metal1 2626 86 2644 90 1 FA0C2
rlabel metal1 2666 46 2684 50 1 FA0C2
rlabel metal1 2754 79 2772 83 1 C0
rlabel metal1 2619 -7 2637 -3 1 FA0S1
rlabel metal1 2661 -7 2679 -3 1 FA0S1not
rlabel metal1 2683 -7 2700 -3 1 FA0S1
rlabel metal1 2700 -131 2718 -127 1 FA0S1
rlabel metal1 2683 -92 2701 -88 1 FA0S1not
rlabel metal1 2699 -46 2717 -42 1 FA0S1not
rlabel metal1 2619 -89 2637 -85 1 D1
rlabel metal1 2661 -89 2679 -85 1 D1not
rlabel metal1 2719 -19 2728 0 1 D1
rlabel metal1 2720 -104 2729 -85 1 D1not
rlabel metal1 2735 -19 2745 36 1 OUT_AS0
rlabel metal1 2736 -104 2745 -49 1 OUT_AS0
rlabel metal1 2469 380 2505 384 5 VDD
rlabel metal1 2469 308 2505 312 1 Gnd
rlabel metal1 2553 329 2562 354 1 D1
rlabel metal1 2554 244 2563 269 1 D1not
rlabel metal1 2453 341 2471 345 1 ASB0
rlabel metal1 2495 341 2513 345 1 ASB0not
rlabel metal1 2533 302 2551 306 1 ASB0not
rlabel metal1 2517 256 2535 260 1 ASB0not
rlabel metal1 2517 341 2534 345 1 ASB0
rlabel metal1 2534 217 2552 221 1 ASB0
rlabel metal1 2570 244 2579 299 1 xorB0
rlabel metal1 2353 344 2389 348 5 VDD
rlabel metal1 2353 272 2389 276 1 Gnd
rlabel metal1 2337 305 2355 309 1 D1
rlabel metal1 2379 305 2397 309 1 D1not
rlabel metal1 2647 380 2683 384 5 VDD
rlabel metal1 2647 308 2683 312 1 Gnd
rlabel metal1 2731 329 2740 354 1 D1
rlabel metal1 2732 244 2741 269 1 D1not
rlabel metal1 2802 380 2838 384 5 VDD
rlabel metal1 2802 308 2838 312 1 Gnd
rlabel metal1 2886 329 2895 354 1 D1
rlabel metal1 2887 244 2896 269 1 D1not
rlabel metal1 2958 380 2994 384 5 VDD
rlabel metal1 2958 308 2994 312 1 Gnd
rlabel metal1 3042 329 3051 354 1 D1
rlabel metal1 3043 244 3052 269 1 D1not
rlabel metal1 2631 341 2649 345 1 ASB1
rlabel metal1 2695 341 2712 345 1 ASB1
rlabel metal1 2712 217 2730 221 1 ASB1
rlabel metal1 2695 256 2713 260 1 ASB1not
rlabel metal1 2711 302 2729 306 1 ASB1not
rlabel metal1 2673 341 2691 345 1 ASB1not
rlabel metal1 2786 341 2804 345 1 ASB2
rlabel metal1 2850 341 2867 345 1 ASB2
rlabel metal1 2867 217 2885 221 1 ASB2
rlabel metal1 2828 341 2846 345 1 ASB2not
rlabel metal1 2866 302 2884 306 1 ASB2not
rlabel metal1 2850 256 2868 260 1 ASB2not
rlabel metal1 2942 341 2960 345 1 ASB3
rlabel metal1 3023 217 3041 221 1 ASB3
rlabel metal1 3006 341 3023 345 1 ASB3
rlabel metal1 3022 302 3040 306 1 ASB3not
rlabel metal1 3006 256 3024 260 1 ASB3not
rlabel metal1 2984 341 3002 345 1 ASB3not
rlabel metal1 3059 244 3068 299 1 xorB3
rlabel metal1 3058 329 3068 384 1 xorB3
rlabel metal1 2902 329 2912 384 1 xorB2
rlabel metal1 2903 244 2912 299 1 xorB2
rlabel metal1 2748 244 2757 299 1 xorB1
rlabel metal1 2747 329 2757 384 1 xorB1
rlabel metal1 2569 329 2579 384 1 xorB0
rlabel metal1 628 -807 776 -803 5 VDD
rlabel metal1 628 -974 776 -970 1 Gnd
rlabel metal1 836 -1012 1040 -1008 1 Gnd
rlabel metal1 836 -806 1040 -802 5 VDD
rlabel metal1 1128 -1012 1332 -1008 1 Gnd
rlabel metal1 1128 -806 1332 -802 5 VDD
rlabel metal1 628 -445 664 -441 5 VDD
rlabel metal1 628 -517 664 -513 1 Gnd
rlabel metal1 628 -527 664 -523 5 VDD
rlabel metal1 628 -599 664 -595 1 Gnd
rlabel metal1 769 -445 805 -441 5 VDD
rlabel metal1 769 -517 805 -513 1 Gnd
rlabel metal1 769 -527 805 -523 5 VDD
rlabel metal1 769 -599 805 -595 1 Gnd
rlabel metal1 628 -626 664 -622 5 VDD
rlabel metal1 628 -698 664 -694 1 Gnd
rlabel metal1 628 -708 664 -704 5 VDD
rlabel metal1 628 -780 664 -776 1 Gnd
rlabel metal1 769 -626 805 -622 5 VDD
rlabel metal1 769 -698 805 -694 1 Gnd
rlabel metal1 769 -708 805 -704 5 VDD
rlabel metal1 769 -780 805 -776 1 Gnd
rlabel metal1 612 -484 630 -480 1 COB0
rlabel metal1 654 -484 672 -480 1 COB0not
rlabel metal1 612 -566 630 -562 1 COA0
rlabel metal1 654 -566 672 -562 1 COA0not
rlabel metal1 753 -484 771 -480 1 COB1
rlabel metal1 795 -484 813 -480 1 COB1not
rlabel metal1 753 -566 771 -562 1 COA1
rlabel metal1 795 -566 813 -562 1 COA1not
rlabel metal1 612 -665 630 -661 1 COB2
rlabel metal1 654 -665 672 -661 1 COB2not
rlabel metal1 612 -747 630 -743 1 COA2
rlabel metal1 654 -747 672 -743 1 COA2not
rlabel metal1 753 -665 771 -661 1 COB3
rlabel metal1 795 -665 813 -661 1 COB3not
rlabel metal1 753 -747 771 -743 1 COA3
rlabel metal1 795 -747 813 -743 1 COA3not
rlabel metal1 675 -484 693 -480 1 COB0
rlabel metal1 692 -523 710 -519 1 COB0not
rlabel metal1 676 -569 694 -565 1 COB0not
rlabel metal1 693 -608 711 -604 1 COB0
rlabel metal1 712 -496 721 -471 1 COA0not
rlabel metal1 713 -581 722 -556 1 COA0
rlabel metal1 728 -496 738 -441 1 EQ1
rlabel metal1 729 -581 738 -526 1 EQ1
rlabel metal1 816 -484 834 -480 1 COB1
rlabel metal1 834 -608 852 -604 1 COB1
rlabel metal1 833 -523 851 -519 1 COB1not
rlabel metal1 817 -569 835 -565 1 COB1not
rlabel metal1 853 -496 862 -471 1 COA1not
rlabel metal1 854 -581 863 -556 1 COA1
rlabel metal1 870 -581 879 -526 1 EQ2
rlabel metal1 869 -496 879 -441 1 EQ2
rlabel metal1 675 -665 693 -661 1 COB2
rlabel metal1 693 -789 711 -785 1 COB2
rlabel metal1 692 -704 710 -700 1 COB2not
rlabel metal1 676 -750 694 -746 1 COB2not
rlabel metal1 713 -762 722 -737 1 COA2
rlabel metal1 712 -677 721 -652 1 COA2not
rlabel metal1 729 -762 738 -707 1 EQ3
rlabel metal1 728 -677 738 -622 1 EQ3
rlabel metal1 869 -677 879 -622 1 EQ4
rlabel metal1 870 -762 879 -707 1 EQ4
rlabel metal1 853 -677 862 -652 1 COA3not
rlabel metal1 854 -762 863 -737 1 COA3
rlabel metal1 816 -665 834 -661 1 COB3
rlabel metal1 834 -789 852 -785 1 COB3
rlabel metal1 833 -704 851 -700 1 COB3not
rlabel metal1 817 -750 835 -746 1 COB3not
rlabel metal1 913 -445 1170 -441 5 VDD
rlabel metal1 913 -651 1170 -647 1 Gnd
rlabel metal1 898 -484 917 -480 1 EQ1
rlabel metal1 926 -500 945 -496 1 EQ1
rlabel metal1 954 -484 973 -480 1 EQ2
rlabel metal1 926 -540 945 -536 1 EQ2
rlabel metal1 1010 -484 1029 -480 1 EQ3
rlabel metal1 926 -580 945 -576 1 EQ3
rlabel metal1 926 -619 945 -615 1 EQ4
rlabel metal1 1066 -484 1085 -480 1 EQ4
rlabel metal1 1158 -493 1177 -489 1 E1
rlabel metal1 943 -790 1035 -786 1 Gnd
rlabel metal1 943 -662 1035 -658 5 VDD
rlabel metal1 1072 -662 1169 -658 5 VDD
rlabel metal1 1072 -794 1169 -790 1 Gnd
rlabel metal1 928 -701 947 -697 1 COA3
rlabel metal1 956 -717 975 -713 1 COA3
rlabel metal1 984 -701 1003 -697 1 COB3not
rlabel metal1 956 -757 975 -753 1 COB3not
rlabel metal1 943 -710 1035 -706 1 G0
rlabel metal1 1083 -701 1101 -697 1 E1
rlabel metal1 1072 -787 1090 -783 1 E1
rlabel metal1 1083 -747 1101 -743 1 G
rlabel metal1 1123 -787 1141 -783 1 G
rlabel metal1 1072 -754 1169 -750 1 L
rlabel metal1 1230 -755 1489 -751 1 Gnd
rlabel metal1 1230 -510 1489 -506 5 VDD
rlabel metal1 669 -846 688 -842 1 COA2
rlabel metal1 641 -902 660 -898 1 COA2
rlabel metal1 725 -846 744 -842 1 COB2not
rlabel metal1 641 -942 660 -938 1 COB2not
rlabel metal1 628 -855 776 -851 1 G1
rlabel metal1 836 -854 1040 -850 1 G2
rlabel metal1 821 -845 840 -841 1 EQ4
rlabel metal1 613 -846 632 -842 1 EQ4
rlabel metal1 641 -862 660 -858 1 EQ4
rlabel metal1 849 -861 868 -857 1 EQ4
rlabel metal1 877 -845 896 -841 1 EQ3
rlabel metal1 849 -901 868 -897 1 EQ3
rlabel metal1 933 -845 952 -841 1 COA1
rlabel metal1 849 -941 868 -937 1 COA1
rlabel metal1 989 -845 1008 -841 1 COB1not
rlabel metal1 849 -980 868 -976 1 COB1not
rlabel metal1 1215 -549 1234 -545 1 EQ4
rlabel metal1 1243 -565 1262 -561 1 EQ4
rlabel metal1 1271 -549 1290 -545 1 EQ3
rlabel metal1 1243 -605 1262 -601 1 EQ3
rlabel metal1 1327 -549 1346 -545 1 EQ2
rlabel metal1 1243 -645 1262 -641 1 EQ2
rlabel metal1 1383 -549 1402 -545 1 COA0
rlabel metal1 1243 -684 1262 -680 1 COA0
rlabel metal1 1438 -549 1457 -545 1 COB0not
rlabel metal1 1243 -723 1262 -719 1 COB0not
rlabel metal1 1230 -558 1489 -554 1 G3
rlabel metal1 1113 -845 1132 -841 1 G0
rlabel metal1 1141 -861 1160 -857 1 G0
rlabel metal1 1169 -845 1188 -841 1 G1
rlabel metal1 1141 -901 1160 -897 1 G1
rlabel metal1 1225 -845 1244 -841 1 G2
rlabel metal1 1141 -941 1160 -937 1 G2
rlabel metal1 1281 -845 1300 -841 1 G3
rlabel metal1 1141 -980 1160 -976 1 G3
rlabel metal1 1128 -854 1332 -850 1 G
rlabel metal1 1410 -1012 1557 -1008 1 Gnd
rlabel metal1 1410 -884 1557 -880 5 VDD
rlabel metal1 1395 -923 1414 -919 1 E1
rlabel metal1 1423 -939 1442 -935 1 E1
rlabel metal1 1451 -923 1470 -919 1 D2
rlabel metal1 1423 -979 1442 -975 1 D2
rlabel metal1 1546 -932 1565 -928 1 E
rlabel metal1 1592 -581 2249 -577 5 VDD
rlabel metal1 1592 -709 2249 -705 1 Gnd
rlabel metal1 1728 -629 1747 -625 1 OUT_AND3
rlabel metal1 1898 -629 1917 -625 1 OUT_AND2
rlabel metal1 2068 -629 2087 -625 1 OUT_AND1
rlabel metal1 2238 -629 2257 -625 1 OUT_AND0
rlabel metal1 1577 -620 1596 -616 1 ANA3
rlabel metal1 1605 -636 1624 -632 1 ANA3
rlabel metal1 1633 -620 1652 -616 1 ANB3
rlabel metal1 1605 -676 1624 -672 1 ANB3
rlabel metal1 1747 -620 1766 -616 1 ANA2
rlabel metal1 1775 -636 1794 -632 1 ANA2
rlabel metal1 1803 -620 1822 -616 1 ANB2
rlabel metal1 1775 -676 1794 -672 1 ANB2
rlabel metal1 1917 -620 1936 -616 1 ANA1
rlabel metal1 1945 -636 1964 -632 1 ANA1
rlabel metal1 1973 -620 1992 -616 1 ANB1
rlabel metal1 1945 -676 1964 -672 1 ANB1
rlabel metal1 2087 -620 2106 -616 1 ANA0
rlabel metal1 2115 -636 2134 -632 1 ANA0
rlabel metal1 2143 -620 2162 -616 1 ANB0
rlabel metal1 2115 -676 2134 -672 1 ANB0
rlabel metal1 993 46 1011 50 1 D0
rlabel metal1 1033 6 1051 10 1 D0
rlabel metal1 1201 239 1220 243 1 A3
rlabel metal1 1376 239 1395 243 1 A2
rlabel metal1 1551 239 1570 243 1 A1
rlabel metal1 1726 239 1745 243 1 A0
rlabel metal1 1698 183 1717 187 1 A0
rlabel metal1 1523 183 1542 187 1 A1
rlabel metal1 1348 183 1367 187 1 A2
rlabel metal1 1173 183 1192 187 1 A3
rlabel metal1 1160 278 1832 282 5 VDD
rlabel metal1 1160 127 1832 131 1 VDD
rlabel metal1 1160 150 1832 154 1 Gnd
rlabel metal1 1201 88 1220 92 1 B3
rlabel metal1 1376 88 1395 92 1 B2
rlabel metal1 1551 88 1570 92 1 B1
rlabel metal1 1726 88 1745 92 1 B0
rlabel metal1 1698 32 1717 36 1 B0
rlabel metal1 1523 32 1542 36 1 B1
rlabel metal1 1348 32 1367 36 1 B2
rlabel metal1 1173 32 1192 36 1 B3
rlabel metal1 1145 239 1164 243 1 DAS
rlabel metal1 1320 239 1339 243 1 DAS
rlabel metal1 1495 239 1514 243 1 DAS
rlabel metal1 1670 239 1689 243 1 DAS
rlabel metal1 1173 223 1192 227 1 DAS
rlabel metal1 1348 223 1367 227 1 DAS
rlabel metal1 1523 223 1542 227 1 DAS
rlabel metal1 1698 223 1717 227 1 DAS
rlabel metal1 1296 230 1315 234 1 ASA3
rlabel metal1 1471 230 1490 234 1 ASA2
rlabel metal1 1646 230 1665 234 1 ASA1
rlabel metal1 1821 230 1840 234 1 ASA0
rlabel metal1 1145 88 1164 92 1 DAS
rlabel metal1 1173 72 1192 76 1 DAS
rlabel metal1 1296 79 1315 83 1 ASB3
rlabel metal1 1320 88 1339 92 1 DAS
rlabel metal1 1348 72 1367 76 1 DAS
rlabel metal1 1471 79 1490 83 1 ASB2
rlabel metal1 1495 88 1514 92 1 DAS
rlabel metal1 1523 72 1542 76 1 DAS
rlabel metal1 1646 79 1665 83 1 ASB1
rlabel metal1 1670 88 1689 92 1 DAS
rlabel metal1 1698 72 1717 76 1 DAS
rlabel metal1 1821 79 1840 83 1 ASB0
rlabel metal1 1160 -1 1840 3 1 Gnd
rlabel metal1 598 541 617 545 1 ANA3
rlabel metal1 773 541 792 545 1 ANA2
rlabel metal1 948 541 967 545 1 ANA1
rlabel metal1 1123 541 1142 545 1 ANA0
rlabel metal1 1123 390 1142 394 1 ANB0
rlabel metal1 948 390 967 394 1 ANB1
rlabel metal1 773 390 792 394 1 ANB2
rlabel metal1 598 390 617 394 1 ANB3
rlabel metal1 475 383 494 387 1 D3
rlabel metal1 447 399 466 403 1 D3
rlabel metal1 650 383 669 387 1 D3
rlabel metal1 622 399 641 403 1 D3
rlabel metal1 825 383 844 387 1 D3
rlabel metal1 797 399 816 403 1 D3
rlabel metal1 1000 383 1019 387 1 D3
rlabel metal1 972 399 991 403 1 D3
rlabel metal1 1000 534 1019 538 1 D3
rlabel metal1 972 550 991 554 1 D3
rlabel metal1 825 534 844 538 1 D3
rlabel metal1 797 550 816 554 1 D3
rlabel metal1 650 534 669 538 1 D3
rlabel metal1 622 550 641 554 1 D3
rlabel metal1 475 534 494 538 1 D3
rlabel metal1 447 550 466 554 1 D3
rlabel metal1 475 343 494 347 1 B3
rlabel metal1 650 343 669 347 1 B2
rlabel metal1 825 343 844 347 1 B1
rlabel metal1 1000 343 1019 347 1 B0
rlabel metal1 1028 399 1047 403 1 B0
rlabel metal1 853 399 872 403 1 B1
rlabel metal1 678 399 697 403 1 B2
rlabel metal1 503 399 522 403 1 B3
rlabel metal1 462 461 1134 465 1 Gnd
rlabel metal1 462 438 1134 442 1 VDD
rlabel metal1 462 589 1134 593 5 VDD
rlabel metal1 475 494 494 498 1 A3
rlabel metal1 650 494 669 498 1 A2
rlabel metal1 825 494 844 498 1 A1
rlabel metal1 1000 494 1019 498 1 A0
rlabel metal1 1028 550 1047 554 1 A0
rlabel metal1 853 550 872 554 1 A1
rlabel metal1 678 550 697 554 1 A2
rlabel metal1 503 550 522 554 1 A3
rlabel metal1 1688 494 1707 498 1 ANB0
rlabel metal1 1716 550 1735 554 1 ANB0
rlabel metal1 1688 534 1707 538 1 ANA0
rlabel metal1 1660 550 1679 554 1 ANA0
rlabel metal1 1518 494 1537 498 1 ANB1
rlabel metal1 1546 550 1565 554 1 ANB1
rlabel metal1 1518 534 1537 538 1 ANA1
rlabel metal1 1490 550 1509 554 1 ANA1
rlabel metal1 1348 494 1367 498 1 ANB2
rlabel metal1 1376 550 1395 554 1 ANB2
rlabel metal1 1348 534 1367 538 1 ANA2
rlabel metal1 1320 550 1339 554 1 ANA2
rlabel metal1 1178 494 1197 498 1 ANB3
rlabel metal1 1206 550 1225 554 1 ANB3
rlabel metal1 1178 534 1197 538 1 ANA3
rlabel metal1 1150 550 1169 554 1 ANA3
rlabel metal1 1811 541 1830 545 1 OUT_AND0
rlabel metal1 1641 541 1660 545 1 OUT_AND1
rlabel metal1 1471 541 1490 545 1 OUT_AND2
rlabel metal1 1301 541 1320 545 1 OUT_AND3
rlabel metal1 1165 461 1822 465 1 Gnd
rlabel metal1 1165 589 1822 593 5 VDD
rlabel metal1 462 310 1142 314 1 Gnd
<< end >>
