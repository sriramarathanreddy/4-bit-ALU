magic
tech scmos
timestamp 1701520416
<< nwell >>
rect 747 401 783 433
rect 803 401 839 433
rect 858 392 894 424
rect 945 401 981 433
rect 1001 401 1037 433
rect 1056 392 1092 424
rect 1137 401 1173 433
rect 1193 401 1229 433
rect 1248 392 1284 424
rect 1339 401 1375 433
rect 1395 401 1431 433
rect 1450 392 1486 424
rect 1542 401 1578 433
rect 1598 401 1634 433
rect 1653 392 1689 424
rect 1745 401 1781 433
rect 1801 401 1837 433
rect 1856 392 1892 424
rect 1949 401 1985 433
rect 2005 401 2041 433
rect 2060 392 2096 424
rect 2152 401 2188 433
rect 2208 401 2244 433
rect 2263 392 2299 424
<< ntransistor >>
rect 790 355 794 375
rect 874 362 878 382
rect 988 355 992 375
rect 1072 362 1076 382
rect 1180 355 1184 375
rect 1264 362 1268 382
rect 1382 355 1386 375
rect 1466 362 1470 382
rect 1585 355 1589 375
rect 1669 362 1673 382
rect 1788 355 1792 375
rect 1872 362 1876 382
rect 1992 355 1996 375
rect 2076 362 2080 382
rect 2195 355 2199 375
rect 2279 362 2283 382
rect 790 315 794 335
rect 988 315 992 335
rect 1180 315 1184 335
rect 1382 315 1386 335
rect 1585 315 1589 335
rect 1788 315 1792 335
rect 1992 315 1996 335
rect 2195 315 2199 335
<< ptransistor >>
rect 764 407 766 427
rect 820 407 822 427
rect 875 398 877 418
rect 962 407 964 427
rect 1018 407 1020 427
rect 1073 398 1075 418
rect 1154 407 1156 427
rect 1210 407 1212 427
rect 1265 398 1267 418
rect 1356 407 1358 427
rect 1412 407 1414 427
rect 1467 398 1469 418
rect 1559 407 1561 427
rect 1615 407 1617 427
rect 1670 398 1672 418
rect 1762 407 1764 427
rect 1818 407 1820 427
rect 1873 398 1875 418
rect 1966 407 1968 427
rect 2022 407 2024 427
rect 2077 398 2079 418
rect 2169 407 2171 427
rect 2225 407 2227 427
rect 2280 398 2282 418
<< ndiffusion >>
rect 789 355 790 375
rect 794 355 795 375
rect 873 362 874 382
rect 878 362 879 382
rect 987 355 988 375
rect 992 355 993 375
rect 1071 362 1072 382
rect 1076 362 1077 382
rect 1179 355 1180 375
rect 1184 355 1185 375
rect 1263 362 1264 382
rect 1268 362 1269 382
rect 1381 355 1382 375
rect 1386 355 1387 375
rect 1465 362 1466 382
rect 1470 362 1471 382
rect 1584 355 1585 375
rect 1589 355 1590 375
rect 1668 362 1669 382
rect 1673 362 1674 382
rect 1787 355 1788 375
rect 1792 355 1793 375
rect 1871 362 1872 382
rect 1876 362 1877 382
rect 1991 355 1992 375
rect 1996 355 1997 375
rect 2075 362 2076 382
rect 2080 362 2081 382
rect 2194 355 2195 375
rect 2199 355 2200 375
rect 2278 362 2279 382
rect 2283 362 2284 382
rect 789 315 790 335
rect 794 315 795 335
rect 987 315 988 335
rect 992 315 993 335
rect 1179 315 1180 335
rect 1184 315 1185 335
rect 1381 315 1382 335
rect 1386 315 1387 335
rect 1584 315 1585 335
rect 1589 315 1590 335
rect 1787 315 1788 335
rect 1792 315 1793 335
rect 1991 315 1992 335
rect 1996 315 1997 335
rect 2194 315 2195 335
rect 2199 315 2200 335
<< pdiffusion >>
rect 763 407 764 427
rect 766 407 767 427
rect 819 407 820 427
rect 822 407 823 427
rect 874 398 875 418
rect 877 398 878 418
rect 961 407 962 427
rect 964 407 965 427
rect 1017 407 1018 427
rect 1020 407 1021 427
rect 1072 398 1073 418
rect 1075 398 1076 418
rect 1153 407 1154 427
rect 1156 407 1157 427
rect 1209 407 1210 427
rect 1212 407 1213 427
rect 1264 398 1265 418
rect 1267 398 1268 418
rect 1355 407 1356 427
rect 1358 407 1359 427
rect 1411 407 1412 427
rect 1414 407 1415 427
rect 1466 398 1467 418
rect 1469 398 1470 418
rect 1558 407 1559 427
rect 1561 407 1562 427
rect 1614 407 1615 427
rect 1617 407 1618 427
rect 1669 398 1670 418
rect 1672 398 1673 418
rect 1761 407 1762 427
rect 1764 407 1765 427
rect 1817 407 1818 427
rect 1820 407 1821 427
rect 1872 398 1873 418
rect 1875 398 1876 418
rect 1965 407 1966 427
rect 1968 407 1969 427
rect 2021 407 2022 427
rect 2024 407 2025 427
rect 2076 398 2077 418
rect 2079 398 2080 418
rect 2168 407 2169 427
rect 2171 407 2172 427
rect 2224 407 2225 427
rect 2227 407 2228 427
rect 2279 398 2280 418
rect 2282 398 2283 418
<< ndcontact >>
rect 779 355 789 375
rect 795 355 805 375
rect 863 362 873 382
rect 879 362 889 382
rect 977 355 987 375
rect 993 355 1003 375
rect 1061 362 1071 382
rect 1077 362 1087 382
rect 1169 355 1179 375
rect 1185 355 1195 375
rect 1253 362 1263 382
rect 1269 362 1279 382
rect 1371 355 1381 375
rect 1387 355 1397 375
rect 1455 362 1465 382
rect 1471 362 1481 382
rect 1574 355 1584 375
rect 1590 355 1600 375
rect 1658 362 1668 382
rect 1674 362 1684 382
rect 1777 355 1787 375
rect 1793 355 1803 375
rect 1861 362 1871 382
rect 1877 362 1887 382
rect 1981 355 1991 375
rect 1997 355 2007 375
rect 2065 362 2075 382
rect 2081 362 2091 382
rect 2184 355 2194 375
rect 2200 355 2210 375
rect 2268 362 2278 382
rect 2284 362 2294 382
rect 779 315 789 335
rect 795 315 805 335
rect 977 315 987 335
rect 993 315 1003 335
rect 1169 315 1179 335
rect 1185 315 1195 335
rect 1371 315 1381 335
rect 1387 315 1397 335
rect 1574 315 1584 335
rect 1590 315 1600 335
rect 1777 315 1787 335
rect 1793 315 1803 335
rect 1981 315 1991 335
rect 1997 315 2007 335
rect 2184 315 2194 335
rect 2200 315 2210 335
<< pdcontact >>
rect 753 407 763 427
rect 767 407 777 427
rect 809 407 819 427
rect 823 407 833 427
rect 864 398 874 418
rect 878 398 888 418
rect 951 407 961 427
rect 965 407 975 427
rect 1007 407 1017 427
rect 1021 407 1031 427
rect 1062 398 1072 418
rect 1076 398 1086 418
rect 1143 407 1153 427
rect 1157 407 1167 427
rect 1199 407 1209 427
rect 1213 407 1223 427
rect 1254 398 1264 418
rect 1268 398 1278 418
rect 1345 407 1355 427
rect 1359 407 1369 427
rect 1401 407 1411 427
rect 1415 407 1425 427
rect 1456 398 1466 418
rect 1470 398 1480 418
rect 1548 407 1558 427
rect 1562 407 1572 427
rect 1604 407 1614 427
rect 1618 407 1628 427
rect 1659 398 1669 418
rect 1673 398 1683 418
rect 1751 407 1761 427
rect 1765 407 1775 427
rect 1807 407 1817 427
rect 1821 407 1831 427
rect 1862 398 1872 418
rect 1876 398 1886 418
rect 1955 407 1965 427
rect 1969 407 1979 427
rect 2011 407 2021 427
rect 2025 407 2035 427
rect 2066 398 2076 418
rect 2080 398 2090 418
rect 2158 407 2168 427
rect 2172 407 2182 427
rect 2214 407 2224 427
rect 2228 407 2238 427
rect 2269 398 2279 418
rect 2283 398 2293 418
<< psubstratepcontact >>
rect 747 305 751 309
rect 835 305 839 309
rect 858 305 862 309
rect 890 305 894 309
rect 945 305 949 309
rect 1033 305 1037 309
rect 1056 305 1060 309
rect 1088 305 1092 309
rect 1137 305 1141 309
rect 1225 305 1229 309
rect 1248 305 1252 309
rect 1280 305 1284 309
rect 1339 305 1343 309
rect 1427 305 1431 309
rect 1450 305 1454 309
rect 1482 305 1486 309
rect 1542 305 1546 309
rect 1630 305 1634 309
rect 1653 305 1657 309
rect 1685 305 1689 309
rect 1745 305 1749 309
rect 1833 305 1837 309
rect 1856 305 1860 309
rect 1888 305 1892 309
rect 1949 305 1953 309
rect 2037 305 2041 309
rect 2060 305 2064 309
rect 2092 305 2096 309
rect 2152 305 2156 309
rect 2240 305 2244 309
rect 2263 305 2267 309
rect 2295 305 2299 309
<< nsubstratencontact >>
rect 747 433 751 437
rect 835 433 839 437
rect 858 433 862 437
rect 890 433 894 437
rect 945 433 949 437
rect 1033 433 1037 437
rect 1056 433 1060 437
rect 1088 433 1092 437
rect 1137 433 1141 437
rect 1225 433 1229 437
rect 1248 433 1252 437
rect 1280 433 1284 437
rect 1339 433 1343 437
rect 1427 433 1431 437
rect 1450 433 1454 437
rect 1482 433 1486 437
rect 1542 433 1546 437
rect 1630 433 1634 437
rect 1653 433 1657 437
rect 1685 433 1689 437
rect 1745 433 1749 437
rect 1833 433 1837 437
rect 1856 433 1860 437
rect 1888 433 1892 437
rect 1949 433 1953 437
rect 2037 433 2041 437
rect 2060 433 2064 437
rect 2092 433 2096 437
rect 2152 433 2156 437
rect 2240 433 2244 437
rect 2263 433 2267 437
rect 2295 433 2299 437
<< polysilicon >>
rect 764 427 766 430
rect 820 427 822 430
rect 875 418 877 421
rect 764 398 766 407
rect 820 398 822 407
rect 930 398 934 440
rect 962 427 964 430
rect 1018 427 1020 430
rect 1073 418 1075 421
rect 962 398 964 407
rect 1018 398 1020 407
rect 1122 398 1126 440
rect 1154 427 1156 430
rect 1210 427 1212 430
rect 1265 418 1267 421
rect 1154 398 1156 407
rect 1210 398 1212 407
rect 1324 398 1328 440
rect 1356 427 1358 430
rect 1412 427 1414 430
rect 1467 418 1469 421
rect 1356 398 1358 407
rect 1412 398 1414 407
rect 1527 398 1531 440
rect 1559 427 1561 430
rect 1615 427 1617 430
rect 1670 418 1672 421
rect 1559 398 1561 407
rect 1615 398 1617 407
rect 1730 398 1734 440
rect 1762 427 1764 430
rect 1818 427 1820 430
rect 1873 418 1875 421
rect 1762 398 1764 407
rect 1818 398 1820 407
rect 1934 398 1938 440
rect 1966 427 1968 430
rect 2022 427 2024 430
rect 2077 418 2079 421
rect 1966 398 1968 407
rect 2022 398 2024 407
rect 2137 398 2141 440
rect 2169 427 2171 430
rect 2225 427 2227 430
rect 2280 418 2282 421
rect 2169 398 2171 407
rect 2225 398 2227 407
rect 751 394 766 398
rect 807 394 822 398
rect 779 378 794 382
rect 790 375 794 378
rect 790 352 794 355
rect 818 342 822 394
rect 875 389 877 398
rect 949 394 964 398
rect 1005 394 1020 398
rect 860 387 877 389
rect 860 385 878 387
rect 874 382 878 385
rect 977 378 992 382
rect 988 375 992 378
rect 874 359 878 362
rect 988 352 992 355
rect 1016 342 1020 394
rect 1073 389 1075 398
rect 1141 394 1156 398
rect 1197 394 1212 398
rect 1058 387 1075 389
rect 1058 385 1076 387
rect 1072 382 1076 385
rect 1169 378 1184 382
rect 1180 375 1184 378
rect 1072 359 1076 362
rect 1180 352 1184 355
rect 1208 342 1212 394
rect 1265 389 1267 398
rect 1343 394 1358 398
rect 1399 394 1414 398
rect 1250 387 1267 389
rect 1250 385 1268 387
rect 1264 382 1268 385
rect 1371 378 1386 382
rect 1382 375 1386 378
rect 1264 359 1268 362
rect 1382 352 1386 355
rect 1410 342 1414 394
rect 1467 389 1469 398
rect 1546 394 1561 398
rect 1602 394 1617 398
rect 1452 387 1469 389
rect 1452 385 1470 387
rect 1466 382 1470 385
rect 1574 378 1589 382
rect 1585 375 1589 378
rect 1466 359 1470 362
rect 1585 352 1589 355
rect 1613 342 1617 394
rect 1670 389 1672 398
rect 1749 394 1764 398
rect 1805 394 1820 398
rect 1655 387 1672 389
rect 1655 385 1673 387
rect 1669 382 1673 385
rect 1777 378 1792 382
rect 1788 375 1792 378
rect 1669 359 1673 362
rect 1788 352 1792 355
rect 1816 342 1820 394
rect 1873 389 1875 398
rect 1953 394 1968 398
rect 2009 394 2024 398
rect 1858 387 1875 389
rect 1858 385 1876 387
rect 1872 382 1876 385
rect 1981 378 1996 382
rect 1992 375 1996 378
rect 1872 359 1876 362
rect 1992 352 1996 355
rect 2020 342 2024 394
rect 2077 389 2079 398
rect 2156 394 2171 398
rect 2212 394 2227 398
rect 2062 387 2079 389
rect 2062 385 2080 387
rect 2076 382 2080 385
rect 2184 378 2199 382
rect 2195 375 2199 378
rect 2076 359 2080 362
rect 2195 352 2199 355
rect 2223 342 2227 394
rect 2280 389 2282 398
rect 2265 387 2282 389
rect 2265 385 2283 387
rect 2279 382 2283 385
rect 2279 359 2283 362
rect 779 338 822 342
rect 977 338 1020 342
rect 1169 338 1212 342
rect 1371 338 1414 342
rect 1574 338 1617 342
rect 1777 338 1820 342
rect 1981 338 2024 342
rect 2184 338 2227 342
rect 790 335 794 338
rect 988 335 992 338
rect 1180 335 1184 338
rect 1382 335 1386 338
rect 1585 335 1589 338
rect 1788 335 1792 338
rect 1992 335 1996 338
rect 2195 335 2199 338
rect 790 312 794 315
rect 988 312 992 315
rect 1180 312 1184 315
rect 1382 312 1386 315
rect 1585 312 1589 315
rect 1788 312 1792 315
rect 1992 312 1996 315
rect 2195 312 2199 315
<< polycontact >>
rect 930 440 934 444
rect 1122 440 1126 444
rect 1324 440 1328 444
rect 1527 440 1531 444
rect 1730 440 1734 444
rect 1934 440 1938 444
rect 2137 440 2141 444
rect 747 394 751 398
rect 775 378 779 382
rect 930 394 934 398
rect 945 394 949 398
rect 856 385 860 389
rect 973 378 977 382
rect 1122 394 1126 398
rect 1137 394 1141 398
rect 1054 385 1058 389
rect 1165 378 1169 382
rect 1324 394 1328 398
rect 1339 394 1343 398
rect 1246 385 1250 389
rect 1367 378 1371 382
rect 1527 394 1531 398
rect 1542 394 1546 398
rect 1448 385 1452 389
rect 1570 378 1574 382
rect 1730 394 1734 398
rect 1745 394 1749 398
rect 1651 385 1655 389
rect 1773 378 1777 382
rect 1934 394 1938 398
rect 1949 394 1953 398
rect 1854 385 1858 389
rect 1977 378 1981 382
rect 2137 394 2141 398
rect 2152 394 2156 398
rect 2058 385 2062 389
rect 2180 378 2184 382
rect 2261 385 2265 389
rect 775 338 779 342
rect 973 338 977 342
rect 1165 338 1169 342
rect 1367 338 1371 342
rect 1570 338 1574 342
rect 1773 338 1777 342
rect 1977 338 1981 342
rect 2180 338 2184 342
<< metal1 >>
rect 732 440 930 444
rect 934 440 1122 444
rect 1126 440 1324 444
rect 1328 440 1527 444
rect 1531 440 1730 444
rect 1734 440 1934 444
rect 1938 440 2137 444
rect 2141 440 2284 444
rect 732 398 736 440
rect 751 433 835 437
rect 839 433 858 437
rect 862 433 890 437
rect 894 433 945 437
rect 949 433 1033 437
rect 1037 433 1056 437
rect 1060 433 1088 437
rect 1092 433 1137 437
rect 1141 433 1225 437
rect 1229 433 1248 437
rect 1252 433 1280 437
rect 1284 433 1339 437
rect 1343 433 1427 437
rect 1431 433 1450 437
rect 1454 433 1482 437
rect 1486 433 1542 437
rect 1546 433 1630 437
rect 1634 433 1653 437
rect 1657 433 1685 437
rect 1689 433 1745 437
rect 1749 433 1833 437
rect 1837 433 1856 437
rect 1860 433 1888 437
rect 1892 433 1949 437
rect 1953 433 2037 437
rect 2041 433 2060 437
rect 2064 433 2092 437
rect 2096 433 2152 437
rect 2156 433 2240 437
rect 2244 433 2263 437
rect 2267 433 2295 437
rect 753 427 763 433
rect 809 427 819 433
rect 732 394 747 398
rect 732 382 736 394
rect 767 389 777 407
rect 823 389 833 407
rect 864 418 874 433
rect 951 427 961 433
rect 1007 427 1017 433
rect 879 389 888 398
rect 934 394 945 398
rect 747 385 856 389
rect 879 385 902 389
rect 732 378 775 382
rect 795 375 805 385
rect 879 382 888 385
rect 930 382 934 394
rect 965 389 975 407
rect 1021 389 1031 407
rect 1062 418 1072 433
rect 1143 427 1153 433
rect 1199 427 1209 433
rect 1077 389 1086 398
rect 1126 394 1137 398
rect 945 385 1054 389
rect 1077 385 1100 389
rect 930 378 973 382
rect 993 375 1003 385
rect 1077 382 1086 385
rect 1122 382 1126 394
rect 1157 389 1167 407
rect 1213 389 1223 407
rect 1254 418 1264 433
rect 1345 427 1355 433
rect 1401 427 1411 433
rect 1269 389 1278 398
rect 1328 394 1339 398
rect 1137 385 1246 389
rect 1269 385 1292 389
rect 779 349 789 355
rect 779 345 805 349
rect 760 338 775 342
rect 795 335 805 345
rect 779 309 789 315
rect 863 309 873 362
rect 1122 378 1165 382
rect 1185 375 1195 385
rect 1269 382 1278 385
rect 1324 382 1328 394
rect 1359 389 1369 407
rect 1415 389 1425 407
rect 1456 418 1466 433
rect 1548 427 1558 433
rect 1604 427 1614 433
rect 1471 389 1480 398
rect 1531 394 1542 398
rect 1339 385 1448 389
rect 1471 385 1494 389
rect 977 349 987 355
rect 977 345 1003 349
rect 958 338 973 342
rect 993 335 1003 345
rect 977 309 987 315
rect 1061 309 1071 362
rect 1324 378 1367 382
rect 1387 375 1397 385
rect 1471 382 1480 385
rect 1527 382 1531 394
rect 1562 389 1572 407
rect 1618 389 1628 407
rect 1659 418 1669 433
rect 1751 427 1761 433
rect 1807 427 1817 433
rect 1674 389 1683 398
rect 1734 394 1745 398
rect 1542 385 1651 389
rect 1674 385 1697 389
rect 1169 349 1179 355
rect 1169 345 1195 349
rect 1150 338 1165 342
rect 1185 335 1195 345
rect 1169 309 1179 315
rect 1253 309 1263 362
rect 1527 378 1570 382
rect 1590 375 1600 385
rect 1674 382 1683 385
rect 1730 382 1734 394
rect 1765 389 1775 407
rect 1821 389 1831 407
rect 1862 418 1872 433
rect 1955 427 1965 433
rect 2011 427 2021 433
rect 1877 389 1886 398
rect 1938 394 1949 398
rect 1745 385 1854 389
rect 1877 385 1900 389
rect 1371 349 1381 355
rect 1371 345 1397 349
rect 1352 338 1367 342
rect 1387 335 1397 345
rect 1371 309 1381 315
rect 1455 309 1465 362
rect 1730 378 1773 382
rect 1793 375 1803 385
rect 1877 382 1886 385
rect 1934 382 1938 394
rect 1969 389 1979 407
rect 2025 389 2035 407
rect 2066 418 2076 433
rect 2158 427 2168 433
rect 2214 427 2224 433
rect 2081 389 2090 398
rect 2141 394 2152 398
rect 1949 385 2058 389
rect 2081 385 2104 389
rect 1574 349 1584 355
rect 1574 345 1600 349
rect 1555 338 1570 342
rect 1590 335 1600 345
rect 1574 309 1584 315
rect 1658 309 1668 362
rect 1934 378 1977 382
rect 1997 375 2007 385
rect 2081 382 2090 385
rect 2137 382 2141 394
rect 2172 389 2182 407
rect 2228 389 2238 407
rect 2269 418 2279 433
rect 2284 389 2293 398
rect 2152 385 2261 389
rect 2284 385 2307 389
rect 1777 349 1787 355
rect 1777 345 1803 349
rect 1758 338 1773 342
rect 1793 335 1803 345
rect 1777 309 1787 315
rect 1861 309 1871 362
rect 2137 378 2180 382
rect 2200 375 2210 385
rect 2284 382 2293 385
rect 1981 349 1991 355
rect 1981 345 2007 349
rect 1962 338 1977 342
rect 1997 335 2007 345
rect 1981 309 1991 315
rect 2065 309 2075 362
rect 2184 349 2194 355
rect 2184 345 2210 349
rect 2165 338 2180 342
rect 2200 335 2210 345
rect 2184 309 2194 315
rect 2268 309 2278 362
rect 751 305 835 309
rect 839 305 858 309
rect 862 305 890 309
rect 894 305 945 309
rect 949 305 1033 309
rect 1037 305 1056 309
rect 1060 305 1088 309
rect 1092 305 1137 309
rect 1141 305 1225 309
rect 1229 305 1248 309
rect 1252 305 1280 309
rect 1284 305 1339 309
rect 1343 305 1427 309
rect 1431 305 1450 309
rect 1454 305 1482 309
rect 1486 305 1542 309
rect 1546 305 1630 309
rect 1634 305 1653 309
rect 1657 305 1685 309
rect 1689 305 1745 309
rect 1749 305 1833 309
rect 1837 305 1856 309
rect 1860 305 1888 309
rect 1892 305 1949 309
rect 1953 305 2037 309
rect 2041 305 2060 309
rect 2064 305 2092 309
rect 2096 305 2152 309
rect 2156 305 2240 309
rect 2244 305 2263 309
rect 2267 305 2295 309
<< labels >>
rlabel metal1 747 433 2299 437 1 VDD
rlabel metal1 747 305 2299 309 1 Gnd
rlabel metal1 732 394 751 398 1 EN
rlabel metal1 760 338 779 342 1 In1
rlabel metal1 958 338 977 342 1 In2
rlabel metal1 1150 338 1169 342 1 In3
rlabel metal1 1352 338 1371 342 1 In4
rlabel metal1 1555 338 1574 342 1 In5
rlabel metal1 1758 338 1777 342 1 In6
rlabel metal1 1962 338 1981 342 1 In7
rlabel metal1 2165 338 2184 342 1 In8
rlabel metal1 888 385 902 389 1 OUT1
rlabel metal1 1086 385 1100 389 1 OUT2
rlabel metal1 1278 385 1292 389 1 OUT3
rlabel metal1 1480 385 1494 389 1 OUT4
rlabel metal1 1683 385 1697 389 1 OUT5
rlabel metal1 1886 385 1900 389 1 OUT6
rlabel metal1 2090 385 2104 389 1 OUT7
rlabel metal1 2293 385 2307 389 1 OUT8
<< end >>
