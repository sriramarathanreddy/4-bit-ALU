magic
tech scmos
timestamp 1701519357
<< nwell >>
rect 236 -102 272 -70
rect 315 -102 351 -70
rect 371 -102 407 -70
rect 426 -111 462 -79
rect 500 -102 536 -70
rect 556 -102 592 -70
rect 611 -111 647 -79
rect 236 -245 272 -213
rect 314 -245 350 -213
rect 370 -245 406 -213
rect 425 -254 461 -222
rect 499 -245 535 -213
rect 555 -245 591 -213
rect 610 -254 646 -222
<< ntransistor >>
rect 252 -188 256 -168
rect 358 -148 362 -128
rect 442 -141 446 -121
rect 543 -148 547 -128
rect 627 -141 631 -121
rect 358 -188 362 -168
rect 543 -188 547 -168
rect 252 -331 256 -311
rect 357 -291 361 -271
rect 441 -284 445 -264
rect 542 -291 546 -271
rect 626 -284 630 -264
rect 357 -331 361 -311
rect 542 -331 546 -311
<< ptransistor >>
rect 253 -96 255 -76
rect 332 -96 334 -76
rect 388 -96 390 -76
rect 443 -105 445 -85
rect 517 -96 519 -76
rect 573 -96 575 -76
rect 628 -105 630 -85
rect 253 -239 255 -219
rect 331 -239 333 -219
rect 387 -239 389 -219
rect 442 -248 444 -228
rect 516 -239 518 -219
rect 572 -239 574 -219
rect 627 -248 629 -228
<< ndiffusion >>
rect 251 -188 252 -168
rect 256 -188 257 -168
rect 357 -148 358 -128
rect 362 -148 363 -128
rect 441 -141 442 -121
rect 446 -141 447 -121
rect 542 -148 543 -128
rect 547 -148 548 -128
rect 626 -141 627 -121
rect 631 -141 632 -121
rect 357 -188 358 -168
rect 362 -188 363 -168
rect 542 -188 543 -168
rect 547 -188 548 -168
rect 251 -331 252 -311
rect 256 -331 257 -311
rect 356 -291 357 -271
rect 361 -291 362 -271
rect 440 -284 441 -264
rect 445 -284 446 -264
rect 541 -291 542 -271
rect 546 -291 547 -271
rect 625 -284 626 -264
rect 630 -284 631 -264
rect 356 -331 357 -311
rect 361 -331 362 -311
rect 541 -331 542 -311
rect 546 -331 547 -311
<< pdiffusion >>
rect 252 -96 253 -76
rect 255 -96 256 -76
rect 331 -96 332 -76
rect 334 -96 335 -76
rect 387 -96 388 -76
rect 390 -96 391 -76
rect 442 -105 443 -85
rect 445 -105 446 -85
rect 516 -96 517 -76
rect 519 -96 520 -76
rect 572 -96 573 -76
rect 575 -96 576 -76
rect 627 -105 628 -85
rect 630 -105 631 -85
rect 252 -239 253 -219
rect 255 -239 256 -219
rect 330 -239 331 -219
rect 333 -239 334 -219
rect 386 -239 387 -219
rect 389 -239 390 -219
rect 441 -248 442 -228
rect 444 -248 445 -228
rect 515 -239 516 -219
rect 518 -239 519 -219
rect 571 -239 572 -219
rect 574 -239 575 -219
rect 626 -248 627 -228
rect 629 -248 630 -228
<< ndcontact >>
rect 241 -188 251 -168
rect 257 -188 267 -168
rect 347 -148 357 -128
rect 363 -148 373 -128
rect 431 -141 441 -121
rect 447 -141 457 -121
rect 532 -148 542 -128
rect 548 -148 558 -128
rect 616 -141 626 -121
rect 632 -141 642 -121
rect 347 -188 357 -168
rect 363 -188 373 -168
rect 532 -188 542 -168
rect 548 -188 558 -168
rect 241 -331 251 -311
rect 257 -331 267 -311
rect 346 -291 356 -271
rect 362 -291 372 -271
rect 430 -284 440 -264
rect 446 -284 456 -264
rect 531 -291 541 -271
rect 547 -291 557 -271
rect 615 -284 625 -264
rect 631 -284 641 -264
rect 346 -331 356 -311
rect 362 -331 372 -311
rect 531 -331 541 -311
rect 547 -331 557 -311
<< pdcontact >>
rect 242 -96 252 -76
rect 256 -96 266 -76
rect 321 -96 331 -76
rect 335 -96 345 -76
rect 377 -96 387 -76
rect 391 -96 401 -76
rect 432 -105 442 -85
rect 446 -105 456 -85
rect 506 -96 516 -76
rect 520 -96 530 -76
rect 562 -96 572 -76
rect 576 -96 586 -76
rect 617 -105 627 -85
rect 631 -105 641 -85
rect 242 -239 252 -219
rect 256 -239 266 -219
rect 320 -239 330 -219
rect 334 -239 344 -219
rect 376 -239 386 -219
rect 390 -239 400 -219
rect 431 -248 441 -228
rect 445 -248 455 -228
rect 505 -239 515 -219
rect 519 -239 529 -219
rect 561 -239 571 -219
rect 575 -239 585 -219
rect 616 -248 626 -228
rect 630 -248 640 -228
<< psubstratepcontact >>
rect 236 -198 240 -194
rect 268 -198 272 -194
rect 315 -198 319 -194
rect 403 -198 407 -194
rect 426 -198 430 -194
rect 458 -198 462 -194
rect 500 -198 504 -194
rect 588 -198 592 -194
rect 611 -198 615 -194
rect 643 -198 647 -194
rect 236 -341 240 -337
rect 268 -341 272 -337
rect 314 -341 318 -337
rect 402 -341 406 -337
rect 425 -341 429 -337
rect 457 -341 461 -337
rect 499 -341 503 -337
rect 587 -341 591 -337
rect 610 -341 614 -337
rect 642 -341 646 -337
<< nsubstratencontact >>
rect 236 -70 240 -66
rect 268 -70 272 -66
rect 315 -70 319 -66
rect 403 -70 407 -66
rect 426 -70 430 -66
rect 458 -70 462 -66
rect 500 -70 504 -66
rect 588 -70 592 -66
rect 611 -70 615 -66
rect 643 -70 647 -66
rect 236 -213 240 -209
rect 268 -213 272 -209
rect 314 -213 318 -209
rect 402 -213 406 -209
rect 425 -213 429 -209
rect 457 -213 461 -209
rect 499 -213 503 -209
rect 587 -213 591 -209
rect 610 -213 614 -209
rect 642 -213 646 -209
<< polysilicon >>
rect 220 -63 480 -59
rect 220 -161 224 -63
rect 253 -76 255 -73
rect 332 -76 334 -73
rect 388 -76 390 -73
rect 443 -85 445 -82
rect 253 -161 255 -96
rect 332 -105 334 -96
rect 388 -105 390 -96
rect 319 -109 334 -105
rect 375 -109 390 -105
rect 347 -125 362 -121
rect 178 -165 220 -161
rect 238 -163 255 -161
rect 238 -165 256 -163
rect 178 -373 182 -165
rect 252 -168 256 -165
rect 252 -191 256 -188
rect 273 -202 277 -165
rect 300 -199 304 -125
rect 358 -128 362 -125
rect 358 -151 362 -148
rect 386 -161 390 -109
rect 443 -114 445 -105
rect 428 -116 445 -114
rect 428 -118 446 -116
rect 442 -121 446 -118
rect 442 -144 446 -141
rect 347 -165 390 -161
rect 475 -161 480 -63
rect 517 -76 519 -73
rect 573 -76 575 -73
rect 628 -85 630 -82
rect 517 -105 519 -96
rect 573 -105 575 -96
rect 504 -109 519 -105
rect 560 -109 575 -105
rect 532 -125 547 -121
rect 543 -128 547 -125
rect 543 -151 547 -148
rect 571 -161 575 -109
rect 628 -114 630 -105
rect 613 -116 630 -114
rect 613 -118 631 -116
rect 627 -121 631 -118
rect 627 -144 631 -141
rect 475 -165 513 -161
rect 532 -165 575 -161
rect 358 -168 362 -165
rect 543 -168 547 -165
rect 358 -191 362 -188
rect 485 -199 489 -185
rect 543 -191 547 -188
rect 211 -206 277 -202
rect 280 -203 513 -199
rect 211 -364 216 -206
rect 253 -219 255 -216
rect 253 -304 255 -239
rect 238 -306 255 -304
rect 280 -304 284 -203
rect 299 -208 488 -206
rect 299 -248 303 -208
rect 331 -219 333 -216
rect 387 -219 389 -216
rect 442 -228 444 -225
rect 331 -248 333 -239
rect 387 -248 389 -239
rect 484 -248 488 -208
rect 516 -219 518 -216
rect 572 -219 574 -216
rect 627 -228 629 -225
rect 516 -248 518 -239
rect 572 -248 574 -239
rect 318 -252 333 -248
rect 374 -252 389 -248
rect 238 -308 256 -306
rect 346 -268 361 -264
rect 220 -344 224 -308
rect 252 -311 256 -308
rect 252 -334 256 -331
rect 299 -344 303 -268
rect 357 -271 361 -268
rect 357 -294 361 -291
rect 385 -304 389 -252
rect 442 -257 444 -248
rect 503 -252 518 -248
rect 559 -252 574 -248
rect 427 -259 444 -257
rect 427 -261 445 -259
rect 441 -264 445 -261
rect 531 -268 546 -264
rect 542 -271 546 -268
rect 441 -287 445 -284
rect 542 -294 546 -291
rect 570 -304 574 -252
rect 627 -257 629 -248
rect 612 -259 629 -257
rect 612 -261 630 -259
rect 626 -264 630 -261
rect 626 -287 630 -284
rect 346 -308 389 -304
rect 531 -308 574 -304
rect 220 -348 303 -344
rect 327 -364 331 -308
rect 357 -311 361 -308
rect 357 -334 361 -331
rect 211 -368 331 -364
rect 512 -373 516 -308
rect 542 -311 546 -308
rect 542 -334 546 -331
rect 178 -377 516 -373
<< polycontact >>
rect 315 -109 319 -105
rect 300 -125 304 -121
rect 343 -125 347 -121
rect 220 -165 224 -161
rect 234 -165 238 -161
rect 273 -165 277 -161
rect 424 -118 428 -114
rect 343 -165 347 -161
rect 500 -109 504 -105
rect 528 -125 532 -121
rect 609 -118 613 -114
rect 513 -165 517 -161
rect 528 -165 532 -161
rect 485 -185 489 -181
rect 220 -308 224 -304
rect 234 -308 238 -304
rect 299 -252 303 -248
rect 314 -252 318 -248
rect 280 -308 284 -304
rect 299 -268 303 -264
rect 342 -268 346 -264
rect 484 -252 488 -248
rect 499 -252 503 -248
rect 423 -261 427 -257
rect 527 -268 531 -264
rect 608 -261 612 -257
rect 327 -308 331 -304
rect 342 -308 346 -304
rect 512 -308 516 -304
rect 527 -308 531 -304
<< metal1 >>
rect 233 -70 236 -66
rect 240 -70 268 -66
rect 272 -70 315 -66
rect 319 -70 403 -66
rect 407 -70 426 -66
rect 430 -70 458 -66
rect 462 -70 500 -66
rect 504 -70 588 -66
rect 592 -70 611 -66
rect 615 -70 643 -66
rect 242 -76 252 -70
rect 321 -76 331 -70
rect 377 -76 387 -70
rect 257 -161 266 -96
rect 300 -109 315 -105
rect 300 -121 304 -109
rect 335 -114 345 -96
rect 391 -114 401 -96
rect 432 -85 442 -70
rect 506 -76 516 -70
rect 562 -76 572 -70
rect 447 -114 456 -105
rect 485 -109 500 -105
rect 315 -118 424 -114
rect 447 -118 470 -114
rect 304 -125 343 -121
rect 363 -128 373 -118
rect 447 -121 456 -118
rect 485 -121 489 -109
rect 520 -114 530 -96
rect 576 -114 586 -96
rect 617 -85 627 -70
rect 632 -114 641 -105
rect 500 -118 609 -114
rect 632 -118 655 -114
rect 485 -125 528 -121
rect 347 -154 357 -148
rect 347 -158 373 -154
rect 224 -165 234 -161
rect 257 -165 273 -161
rect 277 -165 343 -161
rect 257 -168 266 -165
rect 363 -168 373 -158
rect 241 -194 251 -188
rect 347 -194 357 -188
rect 431 -194 441 -141
rect 485 -181 489 -125
rect 548 -128 558 -118
rect 632 -121 641 -118
rect 532 -154 542 -148
rect 532 -158 558 -154
rect 517 -165 528 -161
rect 548 -168 558 -158
rect 532 -194 542 -188
rect 616 -194 626 -141
rect 164 -198 236 -194
rect 240 -198 268 -194
rect 272 -198 315 -194
rect 319 -198 403 -194
rect 407 -198 426 -194
rect 430 -198 458 -194
rect 462 -198 500 -194
rect 504 -198 588 -194
rect 592 -198 611 -194
rect 615 -198 643 -194
rect 164 -337 168 -198
rect 233 -213 236 -209
rect 240 -213 268 -209
rect 272 -213 314 -209
rect 318 -213 402 -209
rect 406 -213 425 -209
rect 429 -213 457 -209
rect 461 -213 499 -209
rect 503 -213 587 -209
rect 591 -213 610 -209
rect 614 -213 642 -209
rect 242 -219 252 -213
rect 320 -219 330 -213
rect 376 -219 386 -213
rect 257 -304 266 -239
rect 303 -252 314 -248
rect 299 -264 303 -252
rect 334 -257 344 -239
rect 390 -257 400 -239
rect 431 -228 441 -213
rect 505 -219 515 -213
rect 561 -219 571 -213
rect 446 -257 455 -248
rect 488 -252 499 -248
rect 314 -261 423 -257
rect 446 -261 469 -257
rect 303 -268 342 -264
rect 362 -271 372 -261
rect 446 -264 455 -261
rect 484 -264 488 -252
rect 519 -257 529 -239
rect 575 -257 585 -239
rect 616 -228 626 -213
rect 631 -257 640 -248
rect 499 -261 608 -257
rect 631 -261 654 -257
rect 484 -268 527 -264
rect 547 -271 557 -261
rect 631 -264 640 -261
rect 346 -297 356 -291
rect 346 -301 372 -297
rect 224 -308 234 -304
rect 257 -308 280 -304
rect 331 -308 342 -304
rect 257 -311 266 -308
rect 362 -311 372 -301
rect 241 -337 251 -331
rect 346 -337 356 -331
rect 430 -337 440 -284
rect 531 -297 541 -291
rect 531 -301 557 -297
rect 516 -308 527 -304
rect 547 -311 557 -301
rect 531 -337 541 -331
rect 615 -337 625 -284
rect 164 -341 236 -337
rect 240 -341 268 -337
rect 272 -341 314 -337
rect 318 -341 402 -337
rect 406 -341 425 -337
rect 429 -341 457 -337
rect 461 -341 499 -337
rect 503 -341 587 -337
rect 591 -341 610 -337
rect 614 -341 642 -337
<< metal2 >>
rect 229 -209 233 -70
<< m123contact >>
rect 228 -70 233 -65
rect 228 -214 233 -209
<< labels >>
rlabel metal1 220 -165 238 -161 1 S0
rlabel metal1 220 -308 238 -304 1 S1
rlabel metal1 266 -165 284 -161 1 S0not
rlabel metal1 266 -308 284 -304 1 S1not
rlabel metal1 456 -118 470 -114 1 D0
rlabel metal1 641 -118 655 -114 1 D1
rlabel metal1 640 -261 654 -257 1 D3
rlabel metal1 455 -261 469 -257 1 D2
rlabel metal1 236 -70 647 -66 1 VDD
rlabel metal1 236 -198 647 -194 1 Gnd
<< end >>
