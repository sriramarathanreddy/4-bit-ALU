module and_4bit_tb;
    reg A3,A2,A1,A0,B3,B2,B0,B1,S1,S0;
    wire OSAC,OSA3,OSA2,OSA1,OSA0,OCl,OCe,OCg,OA3,OA2,OA1,OAS0;

    ALU ALU_tb(/*EN,*/A3,A2,A1,A0,B3,B2,B1,B0,S1,S0,OSAC,OSA3,OSA2,OSA1,OSA0,OCg,OCe,OCl,OA3,OA2,OA1,OAS0);
    initial
    begin
        $dumpfile("ALU_out.vcd");
        $dumpvars(0,ALU_tb);
        $monitor("at T=%4t:A = %b%b%b%b, B = %b%b%b%b,S1 = %b,S0 = %b, Add_Sub = %b%b%b%b%b, is A>B:%b, is A=B:%b, is A<B:%b, AND = %b%b%b%b",$time,A3,A2,A1,A0,B3,B2,B1,B0,S1,S0,OSAC,OSA3,OSA2,OSA1,OSA0,OCg,OCe,OCl,OA3,OA2,OA1,OAS0);
        #2 A3=0;A2=0;A1=0;A0=0;B3=0;B2=0;B1=0;B0=0;S1=0;S0=0;
        #2 A3=0;A2=0;A1=0;A0=0;B3=0;B2=0;B1=0;B0=1;S1=0;S0=0;
        #2 A3=0;A2=0;A1=0;A0=0;B3=0;B2=0;B1=1;B0=0;S1=0;S0=0;
        #2 A3=0;A2=0;A1=0;A0=0;B3=0;B2=0;B1=1;B0=1;S1=0;S0=0;
        #2 A3=0;A2=0;A1=0;A0=0;B3=0;B2=1;B1=0;B0=0;S1=0;S0=0;
        #2 A3=0;A2=0;A1=0;A0=0;B3=0;B2=1;B1=0;B0=1;S1=0;S0=0;
        #2 A3=0;A2=0;A1=0;A0=0;B3=0;B2=1;B1=1;B0=0;S1=0;S0=0;
        #2 A3=0;A2=0;A1=0;A0=0;B3=0;B2=1;B1=1;B0=1;S1=0;S0=0;
        #2 A3=0;A2=0;A1=0;A0=0;B3=1;B2=0;B1=0;B0=0;S1=0;S0=0;
        #2 A3=0;A2=0;A1=0;A0=0;B3=1;B2=0;B1=0;B0=1;S1=0;S0=0;
        #2 A3=0;A2=0;A1=0;A0=0;B3=1;B2=0;B1=1;B0=0;S1=0;S0=0;
        #2 A3=0;A2=0;A1=0;A0=0;B3=1;B2=0;B1=1;B0=1;S1=0;S0=0;
        #2 A3=0;A2=0;A1=0;A0=0;B3=1;B2=1;B1=0;B0=0;S1=0;S0=0;
        #2 A3=0;A2=0;A1=0;A0=0;B3=1;B2=1;B1=0;B0=1;S1=0;S0=0;
        #2 A3=0;A2=0;A1=0;A0=0;B3=1;B2=1;B1=1;B0=0;S1=0;S0=0;
        #2 A3=0;A2=0;A1=0;A0=0;B3=1;B2=1;B1=1;B0=1;S1=0;S0=0;
        #2 A3=0;A2=0;A1=0;A0=1;B3=0;B2=0;B1=0;B0=0;S1=0;S0=0;
        #2 A3=0;A2=0;A1=0;A0=1;B3=0;B2=0;B1=0;B0=1;S1=0;S0=0;
        #2 A3=0;A2=0;A1=0;A0=1;B3=0;B2=0;B1=1;B0=0;S1=0;S0=0;
        #2 A3=0;A2=0;A1=0;A0=1;B3=0;B2=0;B1=1;B0=1;S1=0;S0=0;
        #2 A3=0;A2=0;A1=0;A0=1;B3=0;B2=1;B1=0;B0=0;S1=0;S0=0;
        #2 A3=0;A2=0;A1=0;A0=1;B3=0;B2=1;B1=0;B0=1;S1=0;S0=0;
        #2 A3=0;A2=0;A1=0;A0=1;B3=0;B2=1;B1=1;B0=0;S1=0;S0=0;
        #2 A3=0;A2=0;A1=0;A0=1;B3=0;B2=1;B1=1;B0=1;S1=0;S0=0;
        #2 A3=0;A2=0;A1=0;A0=1;B3=1;B2=0;B1=0;B0=0;S1=0;S0=0;
        #2 A3=0;A2=0;A1=0;A0=1;B3=1;B2=0;B1=0;B0=1;S1=0;S0=0;
        #2 A3=0;A2=0;A1=0;A0=1;B3=1;B2=0;B1=1;B0=0;S1=0;S0=0;
        #2 A3=0;A2=0;A1=0;A0=1;B3=1;B2=0;B1=1;B0=1;S1=0;S0=0;
        #2 A3=0;A2=0;A1=0;A0=1;B3=1;B2=1;B1=0;B0=0;S1=0;S0=0;
        #2 A3=0;A2=0;A1=0;A0=1;B3=1;B2=1;B1=0;B0=1;S1=0;S0=0;
        #2 A3=0;A2=0;A1=0;A0=1;B3=1;B2=1;B1=1;B0=0;S1=0;S0=0;
        #2 A3=0;A2=0;A1=0;A0=1;B3=1;B2=1;B1=1;B0=1;S1=0;S0=0;
        #2 A3=0;A2=0;A1=1;A0=0;B3=0;B2=0;B1=0;B0=0;S1=0;S0=0;
        #2 A3=0;A2=0;A1=1;A0=0;B3=0;B2=0;B1=0;B0=1;S1=0;S0=0;
        #2 A3=0;A2=0;A1=1;A0=0;B3=0;B2=0;B1=1;B0=0;S1=0;S0=0;
        #2 A3=0;A2=0;A1=1;A0=0;B3=0;B2=0;B1=1;B0=1;S1=0;S0=0;
        #2 A3=0;A2=0;A1=1;A0=0;B3=0;B2=1;B1=0;B0=0;S1=0;S0=0;
        #2 A3=0;A2=0;A1=1;A0=0;B3=0;B2=1;B1=0;B0=1;S1=0;S0=0;
        #2 A3=0;A2=0;A1=1;A0=0;B3=0;B2=1;B1=1;B0=0;S1=0;S0=0;
        #2 A3=0;A2=0;A1=1;A0=0;B3=0;B2=1;B1=1;B0=1;S1=0;S0=0;
        #2 A3=0;A2=0;A1=1;A0=0;B3=1;B2=0;B1=0;B0=0;S1=0;S0=0;
        #2 A3=0;A2=0;A1=1;A0=0;B3=1;B2=0;B1=0;B0=1;S1=0;S0=0;
        #2 A3=0;A2=0;A1=1;A0=0;B3=1;B2=0;B1=1;B0=0;S1=0;S0=0;
        #2 A3=0;A2=0;A1=1;A0=0;B3=1;B2=0;B1=1;B0=1;S1=0;S0=0;
        #2 A3=0;A2=0;A1=1;A0=0;B3=1;B2=1;B1=0;B0=0;S1=0;S0=0;
        #2 A3=0;A2=0;A1=1;A0=0;B3=1;B2=1;B1=0;B0=1;S1=0;S0=0;
        #2 A3=0;A2=0;A1=1;A0=0;B3=1;B2=1;B1=1;B0=0;S1=0;S0=0;
        #2 A3=0;A2=0;A1=1;A0=0;B3=1;B2=1;B1=1;B0=1;S1=0;S0=0;
        #2 A3=0;A2=0;A1=1;A0=1;B3=0;B2=0;B1=0;B0=0;S1=0;S0=0;
        #2 A3=0;A2=0;A1=1;A0=1;B3=0;B2=0;B1=0;B0=1;S1=0;S0=0;
        #2 A3=0;A2=0;A1=1;A0=1;B3=0;B2=0;B1=1;B0=0;S1=0;S0=0;
        #2 A3=0;A2=0;A1=1;A0=1;B3=0;B2=0;B1=1;B0=1;S1=0;S0=0;
        #2 A3=0;A2=0;A1=1;A0=1;B3=0;B2=1;B1=0;B0=0;S1=0;S0=0;
        #2 A3=0;A2=0;A1=1;A0=1;B3=0;B2=1;B1=0;B0=1;S1=0;S0=0;
        #2 A3=0;A2=0;A1=1;A0=1;B3=0;B2=1;B1=1;B0=0;S1=0;S0=0;
        #2 A3=0;A2=0;A1=1;A0=1;B3=0;B2=1;B1=1;B0=1;S1=0;S0=0;
        #2 A3=0;A2=0;A1=1;A0=1;B3=1;B2=0;B1=0;B0=0;S1=0;S0=0;
        #2 A3=0;A2=0;A1=1;A0=1;B3=1;B2=0;B1=0;B0=1;S1=0;S0=0;
        #2 A3=0;A2=0;A1=1;A0=1;B3=1;B2=0;B1=1;B0=0;S1=0;S0=0;
        #2 A3=0;A2=0;A1=1;A0=1;B3=1;B2=0;B1=1;B0=1;S1=0;S0=0;
        #2 A3=0;A2=0;A1=1;A0=1;B3=1;B2=1;B1=0;B0=0;S1=0;S0=0;
        #2 A3=0;A2=0;A1=1;A0=1;B3=1;B2=1;B1=0;B0=1;S1=0;S0=0;
        #2 A3=0;A2=0;A1=1;A0=1;B3=1;B2=1;B1=1;B0=0;S1=0;S0=0;
        #2 A3=0;A2=0;A1=1;A0=1;B3=1;B2=1;B1=1;B0=1;S1=0;S0=0;
        #2 A3=0;A2=1;A1=0;A0=0;B3=0;B2=0;B1=0;B0=0;S1=0;S0=0;
        #2 A3=0;A2=1;A1=0;A0=0;B3=0;B2=0;B1=0;B0=1;S1=0;S0=0;
        #2 A3=0;A2=1;A1=0;A0=0;B3=0;B2=0;B1=1;B0=0;S1=0;S0=0;
        #2 A3=0;A2=1;A1=0;A0=0;B3=0;B2=0;B1=1;B0=1;S1=0;S0=0;
        #2 A3=0;A2=1;A1=0;A0=0;B3=0;B2=1;B1=0;B0=0;S1=0;S0=0;
        #2 A3=0;A2=1;A1=0;A0=0;B3=0;B2=1;B1=0;B0=1;S1=0;S0=0;
        #2 A3=0;A2=1;A1=0;A0=0;B3=0;B2=1;B1=1;B0=0;S1=0;S0=0;
        #2 A3=0;A2=1;A1=0;A0=0;B3=0;B2=1;B1=1;B0=1;S1=0;S0=0;
        #2 A3=0;A2=1;A1=0;A0=0;B3=1;B2=0;B1=0;B0=0;S1=0;S0=0;
        #2 A3=0;A2=1;A1=0;A0=0;B3=1;B2=0;B1=0;B0=1;S1=0;S0=0;
        #2 A3=0;A2=1;A1=0;A0=0;B3=1;B2=0;B1=1;B0=0;S1=0;S0=0;
        #2 A3=0;A2=1;A1=0;A0=0;B3=1;B2=0;B1=1;B0=1;S1=0;S0=0;
        #2 A3=0;A2=1;A1=0;A0=0;B3=1;B2=1;B1=0;B0=0;S1=0;S0=0;
        #2 A3=0;A2=1;A1=0;A0=0;B3=1;B2=1;B1=0;B0=1;S1=0;S0=0;
        #2 A3=0;A2=1;A1=0;A0=0;B3=1;B2=1;B1=1;B0=0;S1=0;S0=0;
        #2 A3=0;A2=1;A1=0;A0=0;B3=1;B2=1;B1=1;B0=1;S1=0;S0=0;
        #2 A3=0;A2=1;A1=0;A0=1;B3=0;B2=0;B1=0;B0=0;S1=0;S0=0;
        #2 A3=0;A2=1;A1=0;A0=1;B3=0;B2=0;B1=0;B0=1;S1=0;S0=0;
        #2 A3=0;A2=1;A1=0;A0=1;B3=0;B2=0;B1=1;B0=0;S1=0;S0=0;
        #2 A3=0;A2=1;A1=0;A0=1;B3=0;B2=0;B1=1;B0=1;S1=0;S0=0;
        #2 A3=0;A2=1;A1=0;A0=1;B3=0;B2=1;B1=0;B0=0;S1=0;S0=0;
        #2 A3=0;A2=1;A1=0;A0=1;B3=0;B2=1;B1=0;B0=1;S1=0;S0=0;
        #2 A3=0;A2=1;A1=0;A0=1;B3=0;B2=1;B1=1;B0=0;S1=0;S0=0;
        #2 A3=0;A2=1;A1=0;A0=1;B3=0;B2=1;B1=1;B0=1;S1=0;S0=0;
        #2 A3=0;A2=1;A1=0;A0=1;B3=1;B2=0;B1=0;B0=0;S1=0;S0=0;
        #2 A3=0;A2=1;A1=0;A0=1;B3=1;B2=0;B1=0;B0=1;S1=0;S0=0;
        #2 A3=0;A2=1;A1=0;A0=1;B3=1;B2=0;B1=1;B0=0;S1=0;S0=0;
        #2 A3=0;A2=1;A1=0;A0=1;B3=1;B2=0;B1=1;B0=1;S1=0;S0=0;
        #2 A3=0;A2=1;A1=0;A0=1;B3=1;B2=1;B1=0;B0=0;S1=0;S0=0;
        #2 A3=0;A2=1;A1=0;A0=1;B3=1;B2=1;B1=0;B0=1;S1=0;S0=0;
        #2 A3=0;A2=1;A1=0;A0=1;B3=1;B2=1;B1=1;B0=0;S1=0;S0=0;
        #2 A3=0;A2=1;A1=0;A0=1;B3=1;B2=1;B1=1;B0=1;S1=0;S0=0;
        #2 A3=0;A2=1;A1=1;A0=0;B3=0;B2=0;B1=0;B0=0;S1=0;S0=0;
        #2 A3=0;A2=1;A1=1;A0=0;B3=0;B2=0;B1=0;B0=1;S1=0;S0=0;
        #2 A3=0;A2=1;A1=1;A0=0;B3=0;B2=0;B1=1;B0=0;S1=0;S0=0;
        #2 A3=0;A2=1;A1=1;A0=0;B3=0;B2=0;B1=1;B0=1;S1=0;S0=0;
        #2 A3=0;A2=1;A1=1;A0=0;B3=0;B2=1;B1=0;B0=0;S1=0;S0=0;
        #2 A3=0;A2=1;A1=1;A0=0;B3=0;B2=1;B1=0;B0=1;S1=0;S0=0;
        #2 A3=0;A2=1;A1=1;A0=0;B3=0;B2=1;B1=1;B0=0;S1=0;S0=0;
        #2 A3=0;A2=1;A1=1;A0=0;B3=0;B2=1;B1=1;B0=1;S1=0;S0=0;
        #2 A3=0;A2=1;A1=1;A0=0;B3=1;B2=0;B1=0;B0=0;S1=0;S0=0;
        #2 A3=0;A2=1;A1=1;A0=0;B3=1;B2=0;B1=0;B0=1;S1=0;S0=0;
        #2 A3=0;A2=1;A1=1;A0=0;B3=1;B2=0;B1=1;B0=0;S1=0;S0=0;
        #2 A3=0;A2=1;A1=1;A0=0;B3=1;B2=0;B1=1;B0=1;S1=0;S0=0;
        #2 A3=0;A2=1;A1=1;A0=0;B3=1;B2=1;B1=0;B0=0;S1=0;S0=0;
        #2 A3=0;A2=1;A1=1;A0=0;B3=1;B2=1;B1=0;B0=1;S1=0;S0=0;
        #2 A3=0;A2=1;A1=1;A0=0;B3=1;B2=1;B1=1;B0=0;S1=0;S0=0;
        #2 A3=0;A2=1;A1=1;A0=0;B3=1;B2=1;B1=1;B0=1;S1=0;S0=0;
        #2 A3=0;A2=1;A1=1;A0=1;B3=0;B2=0;B1=0;B0=0;S1=0;S0=0;
        #2 A3=0;A2=1;A1=1;A0=1;B3=0;B2=0;B1=0;B0=1;S1=0;S0=0;
        #2 A3=0;A2=1;A1=1;A0=1;B3=0;B2=0;B1=1;B0=0;S1=0;S0=0;
        #2 A3=0;A2=1;A1=1;A0=1;B3=0;B2=0;B1=1;B0=1;S1=0;S0=0;
        #2 A3=0;A2=1;A1=1;A0=1;B3=0;B2=1;B1=0;B0=0;S1=0;S0=0;
        #2 A3=0;A2=1;A1=1;A0=1;B3=0;B2=1;B1=0;B0=1;S1=0;S0=0;
        #2 A3=0;A2=1;A1=1;A0=1;B3=0;B2=1;B1=1;B0=0;S1=0;S0=0;
        #2 A3=0;A2=1;A1=1;A0=1;B3=0;B2=1;B1=1;B0=1;S1=0;S0=0;
        #2 A3=0;A2=1;A1=1;A0=1;B3=1;B2=0;B1=0;B0=0;S1=0;S0=0;
        #2 A3=0;A2=1;A1=1;A0=1;B3=1;B2=0;B1=0;B0=1;S1=0;S0=0;
        #2 A3=0;A2=1;A1=1;A0=1;B3=1;B2=0;B1=1;B0=0;S1=0;S0=0;
        #2 A3=0;A2=1;A1=1;A0=1;B3=1;B2=0;B1=1;B0=1;S1=0;S0=0;
        #2 A3=0;A2=1;A1=1;A0=1;B3=1;B2=1;B1=0;B0=0;S1=0;S0=0;
        #2 A3=0;A2=1;A1=1;A0=1;B3=1;B2=1;B1=0;B0=1;S1=0;S0=0;
        #2 A3=0;A2=1;A1=1;A0=1;B3=1;B2=1;B1=1;B0=0;S1=0;S0=0;
        #2 A3=0;A2=1;A1=1;A0=1;B3=1;B2=1;B1=1;B0=1;S1=0;S0=0;
        #2 A3=1;A2=0;A1=0;A0=0;B3=0;B2=0;B1=0;B0=0;S1=0;S0=0;
        #2 A3=1;A2=0;A1=0;A0=0;B3=0;B2=0;B1=0;B0=1;S1=0;S0=0;
        #2 A3=1;A2=0;A1=0;A0=0;B3=0;B2=0;B1=1;B0=0;S1=0;S0=0;
        #2 A3=1;A2=0;A1=0;A0=0;B3=0;B2=0;B1=1;B0=1;S1=0;S0=0;
        #2 A3=1;A2=0;A1=0;A0=0;B3=0;B2=1;B1=0;B0=0;S1=0;S0=0;
        #2 A3=1;A2=0;A1=0;A0=0;B3=0;B2=1;B1=0;B0=1;S1=0;S0=0;
        #2 A3=1;A2=0;A1=0;A0=0;B3=0;B2=1;B1=1;B0=0;S1=0;S0=0;
        #2 A3=1;A2=0;A1=0;A0=0;B3=0;B2=1;B1=1;B0=1;S1=0;S0=0;
        #2 A3=1;A2=0;A1=0;A0=0;B3=1;B2=0;B1=0;B0=0;S1=0;S0=0;
        #2 A3=1;A2=0;A1=0;A0=0;B3=1;B2=0;B1=0;B0=1;S1=0;S0=0;
        #2 A3=1;A2=0;A1=0;A0=0;B3=1;B2=0;B1=1;B0=0;S1=0;S0=0;
        #2 A3=1;A2=0;A1=0;A0=0;B3=1;B2=0;B1=1;B0=1;S1=0;S0=0;
        #2 A3=1;A2=0;A1=0;A0=0;B3=1;B2=1;B1=0;B0=0;S1=0;S0=0;
        #2 A3=1;A2=0;A1=0;A0=0;B3=1;B2=1;B1=0;B0=1;S1=0;S0=0;
        #2 A3=1;A2=0;A1=0;A0=0;B3=1;B2=1;B1=1;B0=0;S1=0;S0=0;
        #2 A3=1;A2=0;A1=0;A0=0;B3=1;B2=1;B1=1;B0=1;S1=0;S0=0;
        #2 A3=1;A2=0;A1=0;A0=1;B3=0;B2=0;B1=0;B0=0;S1=0;S0=0;
        #2 A3=1;A2=0;A1=0;A0=1;B3=0;B2=0;B1=0;B0=1;S1=0;S0=0;
        #2 A3=1;A2=0;A1=0;A0=1;B3=0;B2=0;B1=1;B0=0;S1=0;S0=0;
        #2 A3=1;A2=0;A1=0;A0=1;B3=0;B2=0;B1=1;B0=1;S1=0;S0=0;
        #2 A3=1;A2=0;A1=0;A0=1;B3=0;B2=1;B1=0;B0=0;S1=0;S0=0;
        #2 A3=1;A2=0;A1=0;A0=1;B3=0;B2=1;B1=0;B0=1;S1=0;S0=0;
        #2 A3=1;A2=0;A1=0;A0=1;B3=0;B2=1;B1=1;B0=0;S1=0;S0=0;
        #2 A3=1;A2=0;A1=0;A0=1;B3=0;B2=1;B1=1;B0=1;S1=0;S0=0;
        #2 A3=1;A2=0;A1=0;A0=1;B3=1;B2=0;B1=0;B0=0;S1=0;S0=0;
        #2 A3=1;A2=0;A1=0;A0=1;B3=1;B2=0;B1=0;B0=1;S1=0;S0=0;
        #2 A3=1;A2=0;A1=0;A0=1;B3=1;B2=0;B1=1;B0=0;S1=0;S0=0;
        #2 A3=1;A2=0;A1=0;A0=1;B3=1;B2=0;B1=1;B0=1;S1=0;S0=0;
        #2 A3=1;A2=0;A1=0;A0=1;B3=1;B2=1;B1=0;B0=0;S1=0;S0=0;
        #2 A3=1;A2=0;A1=0;A0=1;B3=1;B2=1;B1=0;B0=1;S1=0;S0=0;
        #2 A3=1;A2=0;A1=0;A0=1;B3=1;B2=1;B1=1;B0=0;S1=0;S0=0;
        #2 A3=1;A2=0;A1=0;A0=1;B3=1;B2=1;B1=1;B0=1;S1=0;S0=0;
        #2 A3=1;A2=0;A1=1;A0=0;B3=0;B2=0;B1=0;B0=0;S1=0;S0=0;
        #2 A3=1;A2=0;A1=1;A0=0;B3=0;B2=0;B1=0;B0=1;S1=0;S0=0;
        #2 A3=1;A2=0;A1=1;A0=0;B3=0;B2=0;B1=1;B0=0;S1=0;S0=0;
        #2 A3=1;A2=0;A1=1;A0=0;B3=0;B2=0;B1=1;B0=1;S1=0;S0=0;
        #2 A3=1;A2=0;A1=1;A0=0;B3=0;B2=1;B1=0;B0=0;S1=0;S0=0;
        #2 A3=1;A2=0;A1=1;A0=0;B3=0;B2=1;B1=0;B0=1;S1=0;S0=0;
        #2 A3=1;A2=0;A1=1;A0=0;B3=0;B2=1;B1=1;B0=0;S1=0;S0=0;
        #2 A3=1;A2=0;A1=1;A0=0;B3=0;B2=1;B1=1;B0=1;S1=0;S0=0;
        #2 A3=1;A2=0;A1=1;A0=0;B3=1;B2=0;B1=0;B0=0;S1=0;S0=0;
        #2 A3=1;A2=0;A1=1;A0=0;B3=1;B2=0;B1=0;B0=1;S1=0;S0=0;
        #2 A3=1;A2=0;A1=1;A0=0;B3=1;B2=0;B1=1;B0=0;S1=0;S0=0;
        #2 A3=1;A2=0;A1=1;A0=0;B3=1;B2=0;B1=1;B0=1;S1=0;S0=0;
        #2 A3=1;A2=0;A1=1;A0=0;B3=1;B2=1;B1=0;B0=0;S1=0;S0=0;
        #2 A3=1;A2=0;A1=1;A0=0;B3=1;B2=1;B1=0;B0=1;S1=0;S0=0;
        #2 A3=1;A2=0;A1=1;A0=0;B3=1;B2=1;B1=1;B0=0;S1=0;S0=0;
        #2 A3=1;A2=0;A1=1;A0=0;B3=1;B2=1;B1=1;B0=1;S1=0;S0=0;
        #2 A3=1;A2=0;A1=1;A0=1;B3=0;B2=0;B1=0;B0=0;S1=0;S0=0;
        #2 A3=1;A2=0;A1=1;A0=1;B3=0;B2=0;B1=0;B0=1;S1=0;S0=0;
        #2 A3=1;A2=0;A1=1;A0=1;B3=0;B2=0;B1=1;B0=0;S1=0;S0=0;
        #2 A3=1;A2=0;A1=1;A0=1;B3=0;B2=0;B1=1;B0=1;S1=0;S0=0;
        #2 A3=1;A2=0;A1=1;A0=1;B3=0;B2=1;B1=0;B0=0;S1=0;S0=0;
        #2 A3=1;A2=0;A1=1;A0=1;B3=0;B2=1;B1=0;B0=1;S1=0;S0=0;
        #2 A3=1;A2=0;A1=1;A0=1;B3=0;B2=1;B1=1;B0=0;S1=0;S0=0;
        #2 A3=1;A2=0;A1=1;A0=1;B3=0;B2=1;B1=1;B0=1;S1=0;S0=0;
        #2 A3=1;A2=0;A1=1;A0=1;B3=1;B2=0;B1=0;B0=0;S1=0;S0=0;
        #2 A3=1;A2=0;A1=1;A0=1;B3=1;B2=0;B1=0;B0=1;S1=0;S0=0;
        #2 A3=1;A2=0;A1=1;A0=1;B3=1;B2=0;B1=1;B0=0;S1=0;S0=0;
        #2 A3=1;A2=0;A1=1;A0=1;B3=1;B2=0;B1=1;B0=1;S1=0;S0=0;
        #2 A3=1;A2=0;A1=1;A0=1;B3=1;B2=1;B1=0;B0=0;S1=0;S0=0;
        #2 A3=1;A2=0;A1=1;A0=1;B3=1;B2=1;B1=0;B0=1;S1=0;S0=0;
        #2 A3=1;A2=0;A1=1;A0=1;B3=1;B2=1;B1=1;B0=0;S1=0;S0=0;
        #2 A3=1;A2=0;A1=1;A0=1;B3=1;B2=1;B1=1;B0=1;S1=0;S0=0;
        #2 A3=1;A2=1;A1=0;A0=0;B3=0;B2=0;B1=0;B0=0;S1=0;S0=0;
        #2 A3=1;A2=1;A1=0;A0=0;B3=0;B2=0;B1=0;B0=1;S1=0;S0=0;
        #2 A3=1;A2=1;A1=0;A0=0;B3=0;B2=0;B1=1;B0=0;S1=0;S0=0;
        #2 A3=1;A2=1;A1=0;A0=0;B3=0;B2=0;B1=1;B0=1;S1=0;S0=0;
        #2 A3=1;A2=1;A1=0;A0=0;B3=0;B2=1;B1=0;B0=0;S1=0;S0=0;
        #2 A3=1;A2=1;A1=0;A0=0;B3=0;B2=1;B1=0;B0=1;S1=0;S0=0;
        #2 A3=1;A2=1;A1=0;A0=0;B3=0;B2=1;B1=1;B0=0;S1=0;S0=0;
        #2 A3=1;A2=1;A1=0;A0=0;B3=0;B2=1;B1=1;B0=1;S1=0;S0=0;
        #2 A3=1;A2=1;A1=0;A0=0;B3=1;B2=0;B1=0;B0=0;S1=0;S0=0;
        #2 A3=1;A2=1;A1=0;A0=0;B3=1;B2=0;B1=0;B0=1;S1=0;S0=0;
        #2 A3=1;A2=1;A1=0;A0=0;B3=1;B2=0;B1=1;B0=0;S1=0;S0=0;
        #2 A3=1;A2=1;A1=0;A0=0;B3=1;B2=0;B1=1;B0=1;S1=0;S0=0;
        #2 A3=1;A2=1;A1=0;A0=0;B3=1;B2=1;B1=0;B0=0;S1=0;S0=0;
        #2 A3=1;A2=1;A1=0;A0=0;B3=1;B2=1;B1=0;B0=1;S1=0;S0=0;
        #2 A3=1;A2=1;A1=0;A0=0;B3=1;B2=1;B1=1;B0=0;S1=0;S0=0;
        #2 A3=1;A2=1;A1=0;A0=0;B3=1;B2=1;B1=1;B0=1;S1=0;S0=0;
        #2 A3=1;A2=1;A1=0;A0=1;B3=0;B2=0;B1=0;B0=0;S1=0;S0=0;
        #2 A3=1;A2=1;A1=0;A0=1;B3=0;B2=0;B1=0;B0=1;S1=0;S0=0;
        #2 A3=1;A2=1;A1=0;A0=1;B3=0;B2=0;B1=1;B0=0;S1=0;S0=0;
        #2 A3=1;A2=1;A1=0;A0=1;B3=0;B2=0;B1=1;B0=1;S1=0;S0=0;
        #2 A3=1;A2=1;A1=0;A0=1;B3=0;B2=1;B1=0;B0=0;S1=0;S0=0;
        #2 A3=1;A2=1;A1=0;A0=1;B3=0;B2=1;B1=0;B0=1;S1=0;S0=0;
        #2 A3=1;A2=1;A1=0;A0=1;B3=0;B2=1;B1=1;B0=0;S1=0;S0=0;
        #2 A3=1;A2=1;A1=0;A0=1;B3=0;B2=1;B1=1;B0=1;S1=0;S0=0;
        #2 A3=1;A2=1;A1=0;A0=1;B3=1;B2=0;B1=0;B0=0;S1=0;S0=0;
        #2 A3=1;A2=1;A1=0;A0=1;B3=1;B2=0;B1=0;B0=1;S1=0;S0=0;
        #2 A3=1;A2=1;A1=0;A0=1;B3=1;B2=0;B1=1;B0=0;S1=0;S0=0;
        #2 A3=1;A2=1;A1=0;A0=1;B3=1;B2=0;B1=1;B0=1;S1=0;S0=0;
        #2 A3=1;A2=1;A1=0;A0=1;B3=1;B2=1;B1=0;B0=0;S1=0;S0=0;
        #2 A3=1;A2=1;A1=0;A0=1;B3=1;B2=1;B1=0;B0=1;S1=0;S0=0;
        #2 A3=1;A2=1;A1=0;A0=1;B3=1;B2=1;B1=1;B0=0;S1=0;S0=0;
        #2 A3=1;A2=1;A1=0;A0=1;B3=1;B2=1;B1=1;B0=1;S1=0;S0=0;
        #2 A3=1;A2=1;A1=1;A0=0;B3=0;B2=0;B1=0;B0=0;S1=0;S0=0;
        #2 A3=1;A2=1;A1=1;A0=0;B3=0;B2=0;B1=0;B0=1;S1=0;S0=0;
        #2 A3=1;A2=1;A1=1;A0=0;B3=0;B2=0;B1=1;B0=0;S1=0;S0=0;
        #2 A3=1;A2=1;A1=1;A0=0;B3=0;B2=0;B1=1;B0=1;S1=0;S0=0;
        #2 A3=1;A2=1;A1=1;A0=0;B3=0;B2=1;B1=0;B0=0;S1=0;S0=0;
        #2 A3=1;A2=1;A1=1;A0=0;B3=0;B2=1;B1=0;B0=1;S1=0;S0=0;
        #2 A3=1;A2=1;A1=1;A0=0;B3=0;B2=1;B1=1;B0=0;S1=0;S0=0;
        #2 A3=1;A2=1;A1=1;A0=0;B3=0;B2=1;B1=1;B0=1;S1=0;S0=0;
        #2 A3=1;A2=1;A1=1;A0=0;B3=1;B2=0;B1=0;B0=0;S1=0;S0=0;
        #2 A3=1;A2=1;A1=1;A0=0;B3=1;B2=0;B1=0;B0=1;S1=0;S0=0;
        #2 A3=1;A2=1;A1=1;A0=0;B3=1;B2=0;B1=1;B0=0;S1=0;S0=0;
        #2 A3=1;A2=1;A1=1;A0=0;B3=1;B2=0;B1=1;B0=1;S1=0;S0=0;
        #2 A3=1;A2=1;A1=1;A0=0;B3=1;B2=1;B1=0;B0=0;S1=0;S0=0;
        #2 A3=1;A2=1;A1=1;A0=0;B3=1;B2=1;B1=0;B0=1;S1=0;S0=0;
        #2 A3=1;A2=1;A1=1;A0=0;B3=1;B2=1;B1=1;B0=0;S1=0;S0=0;
        #2 A3=1;A2=1;A1=1;A0=0;B3=1;B2=1;B1=1;B0=1;S1=0;S0=0;
        #2 A3=1;A2=1;A1=1;A0=1;B3=0;B2=0;B1=0;B0=0;S1=0;S0=0;
        #2 A3=1;A2=1;A1=1;A0=1;B3=0;B2=0;B1=0;B0=1;S1=0;S0=0;
        #2 A3=1;A2=1;A1=1;A0=1;B3=0;B2=0;B1=1;B0=0;S1=0;S0=0;
        #2 A3=1;A2=1;A1=1;A0=1;B3=0;B2=0;B1=1;B0=1;S1=0;S0=0;
        #2 A3=1;A2=1;A1=1;A0=1;B3=0;B2=1;B1=0;B0=0;S1=0;S0=0;
        #2 A3=1;A2=1;A1=1;A0=1;B3=0;B2=1;B1=0;B0=1;S1=0;S0=0;
        #2 A3=1;A2=1;A1=1;A0=1;B3=0;B2=1;B1=1;B0=0;S1=0;S0=0;
        #2 A3=1;A2=1;A1=1;A0=1;B3=0;B2=1;B1=1;B0=1;S1=0;S0=0;
        #2 A3=1;A2=1;A1=1;A0=1;B3=1;B2=0;B1=0;B0=0;S1=0;S0=0;
        #2 A3=1;A2=1;A1=1;A0=1;B3=1;B2=0;B1=0;B0=1;S1=0;S0=0;
        #2 A3=1;A2=1;A1=1;A0=1;B3=1;B2=0;B1=1;B0=0;S1=0;S0=0;
        #2 A3=1;A2=1;A1=1;A0=1;B3=1;B2=0;B1=1;B0=1;S1=0;S0=0;
        #2 A3=1;A2=1;A1=1;A0=1;B3=1;B2=1;B1=0;B0=0;S1=0;S0=0;
        #2 A3=1;A2=1;A1=1;A0=1;B3=1;B2=1;B1=0;B0=1;S1=0;S0=0;
        #2 A3=1;A2=1;A1=1;A0=1;B3=1;B2=1;B1=1;B0=0;S1=0;S0=0;
        #2 A3=1;A2=1;A1=1;A0=1;B3=1;B2=1;B1=1;B0=1;S1=0;S0=0;
        #2 A3=0;A2=0;A1=0;A0=0;B3=0;B2=0;B1=0;B0=0;S1=0;S0=1;
        #2 A3=0;A2=0;A1=0;A0=0;B3=0;B2=0;B1=0;B0=1;S1=0;S0=1;
        #2 A3=0;A2=0;A1=0;A0=0;B3=0;B2=0;B1=1;B0=0;S1=0;S0=1;
        #2 A3=0;A2=0;A1=0;A0=0;B3=0;B2=0;B1=1;B0=1;S1=0;S0=1;
        #2 A3=0;A2=0;A1=0;A0=0;B3=0;B2=1;B1=0;B0=0;S1=0;S0=1;
        #2 A3=0;A2=0;A1=0;A0=0;B3=0;B2=1;B1=0;B0=1;S1=0;S0=1;
        #2 A3=0;A2=0;A1=0;A0=0;B3=0;B2=1;B1=1;B0=0;S1=0;S0=1;
        #2 A3=0;A2=0;A1=0;A0=0;B3=0;B2=1;B1=1;B0=1;S1=0;S0=1;
        #2 A3=0;A2=0;A1=0;A0=0;B3=1;B2=0;B1=0;B0=0;S1=0;S0=1;
        #2 A3=0;A2=0;A1=0;A0=0;B3=1;B2=0;B1=0;B0=1;S1=0;S0=1;
        #2 A3=0;A2=0;A1=0;A0=0;B3=1;B2=0;B1=1;B0=0;S1=0;S0=1;
        #2 A3=0;A2=0;A1=0;A0=0;B3=1;B2=0;B1=1;B0=1;S1=0;S0=1;
        #2 A3=0;A2=0;A1=0;A0=0;B3=1;B2=1;B1=0;B0=0;S1=0;S0=1;
        #2 A3=0;A2=0;A1=0;A0=0;B3=1;B2=1;B1=0;B0=1;S1=0;S0=1;
        #2 A3=0;A2=0;A1=0;A0=0;B3=1;B2=1;B1=1;B0=0;S1=0;S0=1;
        #2 A3=0;A2=0;A1=0;A0=0;B3=1;B2=1;B1=1;B0=1;S1=0;S0=1;
        #2 A3=0;A2=0;A1=0;A0=1;B3=0;B2=0;B1=0;B0=0;S1=0;S0=1;
        #2 A3=0;A2=0;A1=0;A0=1;B3=0;B2=0;B1=0;B0=1;S1=0;S0=1;
        #2 A3=0;A2=0;A1=0;A0=1;B3=0;B2=0;B1=1;B0=0;S1=0;S0=1;
        #2 A3=0;A2=0;A1=0;A0=1;B3=0;B2=0;B1=1;B0=1;S1=0;S0=1;
        #2 A3=0;A2=0;A1=0;A0=1;B3=0;B2=1;B1=0;B0=0;S1=0;S0=1;
        #2 A3=0;A2=0;A1=0;A0=1;B3=0;B2=1;B1=0;B0=1;S1=0;S0=1;
        #2 A3=0;A2=0;A1=0;A0=1;B3=0;B2=1;B1=1;B0=0;S1=0;S0=1;
        #2 A3=0;A2=0;A1=0;A0=1;B3=0;B2=1;B1=1;B0=1;S1=0;S0=1;
        #2 A3=0;A2=0;A1=0;A0=1;B3=1;B2=0;B1=0;B0=0;S1=0;S0=1;
        #2 A3=0;A2=0;A1=0;A0=1;B3=1;B2=0;B1=0;B0=1;S1=0;S0=1;
        #2 A3=0;A2=0;A1=0;A0=1;B3=1;B2=0;B1=1;B0=0;S1=0;S0=1;
        #2 A3=0;A2=0;A1=0;A0=1;B3=1;B2=0;B1=1;B0=1;S1=0;S0=1;
        #2 A3=0;A2=0;A1=0;A0=1;B3=1;B2=1;B1=0;B0=0;S1=0;S0=1;
        #2 A3=0;A2=0;A1=0;A0=1;B3=1;B2=1;B1=0;B0=1;S1=0;S0=1;
        #2 A3=0;A2=0;A1=0;A0=1;B3=1;B2=1;B1=1;B0=0;S1=0;S0=1;
        #2 A3=0;A2=0;A1=0;A0=1;B3=1;B2=1;B1=1;B0=1;S1=0;S0=1;
        #2 A3=0;A2=0;A1=1;A0=0;B3=0;B2=0;B1=0;B0=0;S1=0;S0=1;
        #2 A3=0;A2=0;A1=1;A0=0;B3=0;B2=0;B1=0;B0=1;S1=0;S0=1;
        #2 A3=0;A2=0;A1=1;A0=0;B3=0;B2=0;B1=1;B0=0;S1=0;S0=1;
        #2 A3=0;A2=0;A1=1;A0=0;B3=0;B2=0;B1=1;B0=1;S1=0;S0=1;
        #2 A3=0;A2=0;A1=1;A0=0;B3=0;B2=1;B1=0;B0=0;S1=0;S0=1;
        #2 A3=0;A2=0;A1=1;A0=0;B3=0;B2=1;B1=0;B0=1;S1=0;S0=1;
        #2 A3=0;A2=0;A1=1;A0=0;B3=0;B2=1;B1=1;B0=0;S1=0;S0=1;
        #2 A3=0;A2=0;A1=1;A0=0;B3=0;B2=1;B1=1;B0=1;S1=0;S0=1;
        #2 A3=0;A2=0;A1=1;A0=0;B3=1;B2=0;B1=0;B0=0;S1=0;S0=1;
        #2 A3=0;A2=0;A1=1;A0=0;B3=1;B2=0;B1=0;B0=1;S1=0;S0=1;
        #2 A3=0;A2=0;A1=1;A0=0;B3=1;B2=0;B1=1;B0=0;S1=0;S0=1;
        #2 A3=0;A2=0;A1=1;A0=0;B3=1;B2=0;B1=1;B0=1;S1=0;S0=1;
        #2 A3=0;A2=0;A1=1;A0=0;B3=1;B2=1;B1=0;B0=0;S1=0;S0=1;
        #2 A3=0;A2=0;A1=1;A0=0;B3=1;B2=1;B1=0;B0=1;S1=0;S0=1;
        #2 A3=0;A2=0;A1=1;A0=0;B3=1;B2=1;B1=1;B0=0;S1=0;S0=1;
        #2 A3=0;A2=0;A1=1;A0=0;B3=1;B2=1;B1=1;B0=1;S1=0;S0=1;
        #2 A3=0;A2=0;A1=1;A0=1;B3=0;B2=0;B1=0;B0=0;S1=0;S0=1;
        #2 A3=0;A2=0;A1=1;A0=1;B3=0;B2=0;B1=0;B0=1;S1=0;S0=1;
        #2 A3=0;A2=0;A1=1;A0=1;B3=0;B2=0;B1=1;B0=0;S1=0;S0=1;
        #2 A3=0;A2=0;A1=1;A0=1;B3=0;B2=0;B1=1;B0=1;S1=0;S0=1;
        #2 A3=0;A2=0;A1=1;A0=1;B3=0;B2=1;B1=0;B0=0;S1=0;S0=1;
        #2 A3=0;A2=0;A1=1;A0=1;B3=0;B2=1;B1=0;B0=1;S1=0;S0=1;
        #2 A3=0;A2=0;A1=1;A0=1;B3=0;B2=1;B1=1;B0=0;S1=0;S0=1;
        #2 A3=0;A2=0;A1=1;A0=1;B3=0;B2=1;B1=1;B0=1;S1=0;S0=1;
        #2 A3=0;A2=0;A1=1;A0=1;B3=1;B2=0;B1=0;B0=0;S1=0;S0=1;
        #2 A3=0;A2=0;A1=1;A0=1;B3=1;B2=0;B1=0;B0=1;S1=0;S0=1;
        #2 A3=0;A2=0;A1=1;A0=1;B3=1;B2=0;B1=1;B0=0;S1=0;S0=1;
        #2 A3=0;A2=0;A1=1;A0=1;B3=1;B2=0;B1=1;B0=1;S1=0;S0=1;
        #2 A3=0;A2=0;A1=1;A0=1;B3=1;B2=1;B1=0;B0=0;S1=0;S0=1;
        #2 A3=0;A2=0;A1=1;A0=1;B3=1;B2=1;B1=0;B0=1;S1=0;S0=1;
        #2 A3=0;A2=0;A1=1;A0=1;B3=1;B2=1;B1=1;B0=0;S1=0;S0=1;
        #2 A3=0;A2=0;A1=1;A0=1;B3=1;B2=1;B1=1;B0=1;S1=0;S0=1;
        #2 A3=0;A2=1;A1=0;A0=0;B3=0;B2=0;B1=0;B0=0;S1=0;S0=1;
        #2 A3=0;A2=1;A1=0;A0=0;B3=0;B2=0;B1=0;B0=1;S1=0;S0=1;
        #2 A3=0;A2=1;A1=0;A0=0;B3=0;B2=0;B1=1;B0=0;S1=0;S0=1;
        #2 A3=0;A2=1;A1=0;A0=0;B3=0;B2=0;B1=1;B0=1;S1=0;S0=1;
        #2 A3=0;A2=1;A1=0;A0=0;B3=0;B2=1;B1=0;B0=0;S1=0;S0=1;
        #2 A3=0;A2=1;A1=0;A0=0;B3=0;B2=1;B1=0;B0=1;S1=0;S0=1;
        #2 A3=0;A2=1;A1=0;A0=0;B3=0;B2=1;B1=1;B0=0;S1=0;S0=1;
        #2 A3=0;A2=1;A1=0;A0=0;B3=0;B2=1;B1=1;B0=1;S1=0;S0=1;
        #2 A3=0;A2=1;A1=0;A0=0;B3=1;B2=0;B1=0;B0=0;S1=0;S0=1;
        #2 A3=0;A2=1;A1=0;A0=0;B3=1;B2=0;B1=0;B0=1;S1=0;S0=1;
        #2 A3=0;A2=1;A1=0;A0=0;B3=1;B2=0;B1=1;B0=0;S1=0;S0=1;
        #2 A3=0;A2=1;A1=0;A0=0;B3=1;B2=0;B1=1;B0=1;S1=0;S0=1;
        #2 A3=0;A2=1;A1=0;A0=0;B3=1;B2=1;B1=0;B0=0;S1=0;S0=1;
        #2 A3=0;A2=1;A1=0;A0=0;B3=1;B2=1;B1=0;B0=1;S1=0;S0=1;
        #2 A3=0;A2=1;A1=0;A0=0;B3=1;B2=1;B1=1;B0=0;S1=0;S0=1;
        #2 A3=0;A2=1;A1=0;A0=0;B3=1;B2=1;B1=1;B0=1;S1=0;S0=1;
        #2 A3=0;A2=1;A1=0;A0=1;B3=0;B2=0;B1=0;B0=0;S1=0;S0=1;
        #2 A3=0;A2=1;A1=0;A0=1;B3=0;B2=0;B1=0;B0=1;S1=0;S0=1;
        #2 A3=0;A2=1;A1=0;A0=1;B3=0;B2=0;B1=1;B0=0;S1=0;S0=1;
        #2 A3=0;A2=1;A1=0;A0=1;B3=0;B2=0;B1=1;B0=1;S1=0;S0=1;
        #2 A3=0;A2=1;A1=0;A0=1;B3=0;B2=1;B1=0;B0=0;S1=0;S0=1;
        #2 A3=0;A2=1;A1=0;A0=1;B3=0;B2=1;B1=0;B0=1;S1=0;S0=1;
        #2 A3=0;A2=1;A1=0;A0=1;B3=0;B2=1;B1=1;B0=0;S1=0;S0=1;
        #2 A3=0;A2=1;A1=0;A0=1;B3=0;B2=1;B1=1;B0=1;S1=0;S0=1;
        #2 A3=0;A2=1;A1=0;A0=1;B3=1;B2=0;B1=0;B0=0;S1=0;S0=1;
        #2 A3=0;A2=1;A1=0;A0=1;B3=1;B2=0;B1=0;B0=1;S1=0;S0=1;
        #2 A3=0;A2=1;A1=0;A0=1;B3=1;B2=0;B1=1;B0=0;S1=0;S0=1;
        #2 A3=0;A2=1;A1=0;A0=1;B3=1;B2=0;B1=1;B0=1;S1=0;S0=1;
        #2 A3=0;A2=1;A1=0;A0=1;B3=1;B2=1;B1=0;B0=0;S1=0;S0=1;
        #2 A3=0;A2=1;A1=0;A0=1;B3=1;B2=1;B1=0;B0=1;S1=0;S0=1;
        #2 A3=0;A2=1;A1=0;A0=1;B3=1;B2=1;B1=1;B0=0;S1=0;S0=1;
        #2 A3=0;A2=1;A1=0;A0=1;B3=1;B2=1;B1=1;B0=1;S1=0;S0=1;
        #2 A3=0;A2=1;A1=1;A0=0;B3=0;B2=0;B1=0;B0=0;S1=0;S0=1;
        #2 A3=0;A2=1;A1=1;A0=0;B3=0;B2=0;B1=0;B0=1;S1=0;S0=1;
        #2 A3=0;A2=1;A1=1;A0=0;B3=0;B2=0;B1=1;B0=0;S1=0;S0=1;
        #2 A3=0;A2=1;A1=1;A0=0;B3=0;B2=0;B1=1;B0=1;S1=0;S0=1;
        #2 A3=0;A2=1;A1=1;A0=0;B3=0;B2=1;B1=0;B0=0;S1=0;S0=1;
        #2 A3=0;A2=1;A1=1;A0=0;B3=0;B2=1;B1=0;B0=1;S1=0;S0=1;
        #2 A3=0;A2=1;A1=1;A0=0;B3=0;B2=1;B1=1;B0=0;S1=0;S0=1;
        #2 A3=0;A2=1;A1=1;A0=0;B3=0;B2=1;B1=1;B0=1;S1=0;S0=1;
        #2 A3=0;A2=1;A1=1;A0=0;B3=1;B2=0;B1=0;B0=0;S1=0;S0=1;
        #2 A3=0;A2=1;A1=1;A0=0;B3=1;B2=0;B1=0;B0=1;S1=0;S0=1;
        #2 A3=0;A2=1;A1=1;A0=0;B3=1;B2=0;B1=1;B0=0;S1=0;S0=1;
        #2 A3=0;A2=1;A1=1;A0=0;B3=1;B2=0;B1=1;B0=1;S1=0;S0=1;
        #2 A3=0;A2=1;A1=1;A0=0;B3=1;B2=1;B1=0;B0=0;S1=0;S0=1;
        #2 A3=0;A2=1;A1=1;A0=0;B3=1;B2=1;B1=0;B0=1;S1=0;S0=1;
        #2 A3=0;A2=1;A1=1;A0=0;B3=1;B2=1;B1=1;B0=0;S1=0;S0=1;
        #2 A3=0;A2=1;A1=1;A0=0;B3=1;B2=1;B1=1;B0=1;S1=0;S0=1;
        #2 A3=0;A2=1;A1=1;A0=1;B3=0;B2=0;B1=0;B0=0;S1=0;S0=1;
        #2 A3=0;A2=1;A1=1;A0=1;B3=0;B2=0;B1=0;B0=1;S1=0;S0=1;
        #2 A3=0;A2=1;A1=1;A0=1;B3=0;B2=0;B1=1;B0=0;S1=0;S0=1;
        #2 A3=0;A2=1;A1=1;A0=1;B3=0;B2=0;B1=1;B0=1;S1=0;S0=1;
        #2 A3=0;A2=1;A1=1;A0=1;B3=0;B2=1;B1=0;B0=0;S1=0;S0=1;
        #2 A3=0;A2=1;A1=1;A0=1;B3=0;B2=1;B1=0;B0=1;S1=0;S0=1;
        #2 A3=0;A2=1;A1=1;A0=1;B3=0;B2=1;B1=1;B0=0;S1=0;S0=1;
        #2 A3=0;A2=1;A1=1;A0=1;B3=0;B2=1;B1=1;B0=1;S1=0;S0=1;
        #2 A3=0;A2=1;A1=1;A0=1;B3=1;B2=0;B1=0;B0=0;S1=0;S0=1;
        #2 A3=0;A2=1;A1=1;A0=1;B3=1;B2=0;B1=0;B0=1;S1=0;S0=1;
        #2 A3=0;A2=1;A1=1;A0=1;B3=1;B2=0;B1=1;B0=0;S1=0;S0=1;
        #2 A3=0;A2=1;A1=1;A0=1;B3=1;B2=0;B1=1;B0=1;S1=0;S0=1;
        #2 A3=0;A2=1;A1=1;A0=1;B3=1;B2=1;B1=0;B0=0;S1=0;S0=1;
        #2 A3=0;A2=1;A1=1;A0=1;B3=1;B2=1;B1=0;B0=1;S1=0;S0=1;
        #2 A3=0;A2=1;A1=1;A0=1;B3=1;B2=1;B1=1;B0=0;S1=0;S0=1;
        #2 A3=0;A2=1;A1=1;A0=1;B3=1;B2=1;B1=1;B0=1;S1=0;S0=1;
        #2 A3=1;A2=0;A1=0;A0=0;B3=0;B2=0;B1=0;B0=0;S1=0;S0=1;
        #2 A3=1;A2=0;A1=0;A0=0;B3=0;B2=0;B1=0;B0=1;S1=0;S0=1;
        #2 A3=1;A2=0;A1=0;A0=0;B3=0;B2=0;B1=1;B0=0;S1=0;S0=1;
        #2 A3=1;A2=0;A1=0;A0=0;B3=0;B2=0;B1=1;B0=1;S1=0;S0=1;
        #2 A3=1;A2=0;A1=0;A0=0;B3=0;B2=1;B1=0;B0=0;S1=0;S0=1;
        #2 A3=1;A2=0;A1=0;A0=0;B3=0;B2=1;B1=0;B0=1;S1=0;S0=1;
        #2 A3=1;A2=0;A1=0;A0=0;B3=0;B2=1;B1=1;B0=0;S1=0;S0=1;
        #2 A3=1;A2=0;A1=0;A0=0;B3=0;B2=1;B1=1;B0=1;S1=0;S0=1;
        #2 A3=1;A2=0;A1=0;A0=0;B3=1;B2=0;B1=0;B0=0;S1=0;S0=1;
        #2 A3=1;A2=0;A1=0;A0=0;B3=1;B2=0;B1=0;B0=1;S1=0;S0=1;
        #2 A3=1;A2=0;A1=0;A0=0;B3=1;B2=0;B1=1;B0=0;S1=0;S0=1;
        #2 A3=1;A2=0;A1=0;A0=0;B3=1;B2=0;B1=1;B0=1;S1=0;S0=1;
        #2 A3=1;A2=0;A1=0;A0=0;B3=1;B2=1;B1=0;B0=0;S1=0;S0=1;
        #2 A3=1;A2=0;A1=0;A0=0;B3=1;B2=1;B1=0;B0=1;S1=0;S0=1;
        #2 A3=1;A2=0;A1=0;A0=0;B3=1;B2=1;B1=1;B0=0;S1=0;S0=1;
        #2 A3=1;A2=0;A1=0;A0=0;B3=1;B2=1;B1=1;B0=1;S1=0;S0=1;
        #2 A3=1;A2=0;A1=0;A0=1;B3=0;B2=0;B1=0;B0=0;S1=0;S0=1;
        #2 A3=1;A2=0;A1=0;A0=1;B3=0;B2=0;B1=0;B0=1;S1=0;S0=1;
        #2 A3=1;A2=0;A1=0;A0=1;B3=0;B2=0;B1=1;B0=0;S1=0;S0=1;
        #2 A3=1;A2=0;A1=0;A0=1;B3=0;B2=0;B1=1;B0=1;S1=0;S0=1;
        #2 A3=1;A2=0;A1=0;A0=1;B3=0;B2=1;B1=0;B0=0;S1=0;S0=1;
        #2 A3=1;A2=0;A1=0;A0=1;B3=0;B2=1;B1=0;B0=1;S1=0;S0=1;
        #2 A3=1;A2=0;A1=0;A0=1;B3=0;B2=1;B1=1;B0=0;S1=0;S0=1;
        #2 A3=1;A2=0;A1=0;A0=1;B3=0;B2=1;B1=1;B0=1;S1=0;S0=1;
        #2 A3=1;A2=0;A1=0;A0=1;B3=1;B2=0;B1=0;B0=0;S1=0;S0=1;
        #2 A3=1;A2=0;A1=0;A0=1;B3=1;B2=0;B1=0;B0=1;S1=0;S0=1;
        #2 A3=1;A2=0;A1=0;A0=1;B3=1;B2=0;B1=1;B0=0;S1=0;S0=1;
        #2 A3=1;A2=0;A1=0;A0=1;B3=1;B2=0;B1=1;B0=1;S1=0;S0=1;
        #2 A3=1;A2=0;A1=0;A0=1;B3=1;B2=1;B1=0;B0=0;S1=0;S0=1;
        #2 A3=1;A2=0;A1=0;A0=1;B3=1;B2=1;B1=0;B0=1;S1=0;S0=1;
        #2 A3=1;A2=0;A1=0;A0=1;B3=1;B2=1;B1=1;B0=0;S1=0;S0=1;
        #2 A3=1;A2=0;A1=0;A0=1;B3=1;B2=1;B1=1;B0=1;S1=0;S0=1;
        #2 A3=1;A2=0;A1=1;A0=0;B3=0;B2=0;B1=0;B0=0;S1=0;S0=1;
        #2 A3=1;A2=0;A1=1;A0=0;B3=0;B2=0;B1=0;B0=1;S1=0;S0=1;
        #2 A3=1;A2=0;A1=1;A0=0;B3=0;B2=0;B1=1;B0=0;S1=0;S0=1;
        #2 A3=1;A2=0;A1=1;A0=0;B3=0;B2=0;B1=1;B0=1;S1=0;S0=1;
        #2 A3=1;A2=0;A1=1;A0=0;B3=0;B2=1;B1=0;B0=0;S1=0;S0=1;
        #2 A3=1;A2=0;A1=1;A0=0;B3=0;B2=1;B1=0;B0=1;S1=0;S0=1;
        #2 A3=1;A2=0;A1=1;A0=0;B3=0;B2=1;B1=1;B0=0;S1=0;S0=1;
        #2 A3=1;A2=0;A1=1;A0=0;B3=0;B2=1;B1=1;B0=1;S1=0;S0=1;
        #2 A3=1;A2=0;A1=1;A0=0;B3=1;B2=0;B1=0;B0=0;S1=0;S0=1;
        #2 A3=1;A2=0;A1=1;A0=0;B3=1;B2=0;B1=0;B0=1;S1=0;S0=1;
        #2 A3=1;A2=0;A1=1;A0=0;B3=1;B2=0;B1=1;B0=0;S1=0;S0=1;
        #2 A3=1;A2=0;A1=1;A0=0;B3=1;B2=0;B1=1;B0=1;S1=0;S0=1;
        #2 A3=1;A2=0;A1=1;A0=0;B3=1;B2=1;B1=0;B0=0;S1=0;S0=1;
        #2 A3=1;A2=0;A1=1;A0=0;B3=1;B2=1;B1=0;B0=1;S1=0;S0=1;
        #2 A3=1;A2=0;A1=1;A0=0;B3=1;B2=1;B1=1;B0=0;S1=0;S0=1;
        #2 A3=1;A2=0;A1=1;A0=0;B3=1;B2=1;B1=1;B0=1;S1=0;S0=1;
        #2 A3=1;A2=0;A1=1;A0=1;B3=0;B2=0;B1=0;B0=0;S1=0;S0=1;
        #2 A3=1;A2=0;A1=1;A0=1;B3=0;B2=0;B1=0;B0=1;S1=0;S0=1;
        #2 A3=1;A2=0;A1=1;A0=1;B3=0;B2=0;B1=1;B0=0;S1=0;S0=1;
        #2 A3=1;A2=0;A1=1;A0=1;B3=0;B2=0;B1=1;B0=1;S1=0;S0=1;
        #2 A3=1;A2=0;A1=1;A0=1;B3=0;B2=1;B1=0;B0=0;S1=0;S0=1;
        #2 A3=1;A2=0;A1=1;A0=1;B3=0;B2=1;B1=0;B0=1;S1=0;S0=1;
        #2 A3=1;A2=0;A1=1;A0=1;B3=0;B2=1;B1=1;B0=0;S1=0;S0=1;
        #2 A3=1;A2=0;A1=1;A0=1;B3=0;B2=1;B1=1;B0=1;S1=0;S0=1;
        #2 A3=1;A2=0;A1=1;A0=1;B3=1;B2=0;B1=0;B0=0;S1=0;S0=1;
        #2 A3=1;A2=0;A1=1;A0=1;B3=1;B2=0;B1=0;B0=1;S1=0;S0=1;
        #2 A3=1;A2=0;A1=1;A0=1;B3=1;B2=0;B1=1;B0=0;S1=0;S0=1;
        #2 A3=1;A2=0;A1=1;A0=1;B3=1;B2=0;B1=1;B0=1;S1=0;S0=1;
        #2 A3=1;A2=0;A1=1;A0=1;B3=1;B2=1;B1=0;B0=0;S1=0;S0=1;
        #2 A3=1;A2=0;A1=1;A0=1;B3=1;B2=1;B1=0;B0=1;S1=0;S0=1;
        #2 A3=1;A2=0;A1=1;A0=1;B3=1;B2=1;B1=1;B0=0;S1=0;S0=1;
        #2 A3=1;A2=0;A1=1;A0=1;B3=1;B2=1;B1=1;B0=1;S1=0;S0=1;
        #2 A3=1;A2=1;A1=0;A0=0;B3=0;B2=0;B1=0;B0=0;S1=0;S0=1;
        #2 A3=1;A2=1;A1=0;A0=0;B3=0;B2=0;B1=0;B0=1;S1=0;S0=1;
        #2 A3=1;A2=1;A1=0;A0=0;B3=0;B2=0;B1=1;B0=0;S1=0;S0=1;
        #2 A3=1;A2=1;A1=0;A0=0;B3=0;B2=0;B1=1;B0=1;S1=0;S0=1;
        #2 A3=1;A2=1;A1=0;A0=0;B3=0;B2=1;B1=0;B0=0;S1=0;S0=1;
        #2 A3=1;A2=1;A1=0;A0=0;B3=0;B2=1;B1=0;B0=1;S1=0;S0=1;
        #2 A3=1;A2=1;A1=0;A0=0;B3=0;B2=1;B1=1;B0=0;S1=0;S0=1;
        #2 A3=1;A2=1;A1=0;A0=0;B3=0;B2=1;B1=1;B0=1;S1=0;S0=1;
        #2 A3=1;A2=1;A1=0;A0=0;B3=1;B2=0;B1=0;B0=0;S1=0;S0=1;
        #2 A3=1;A2=1;A1=0;A0=0;B3=1;B2=0;B1=0;B0=1;S1=0;S0=1;
        #2 A3=1;A2=1;A1=0;A0=0;B3=1;B2=0;B1=1;B0=0;S1=0;S0=1;
        #2 A3=1;A2=1;A1=0;A0=0;B3=1;B2=0;B1=1;B0=1;S1=0;S0=1;
        #2 A3=1;A2=1;A1=0;A0=0;B3=1;B2=1;B1=0;B0=0;S1=0;S0=1;
        #2 A3=1;A2=1;A1=0;A0=0;B3=1;B2=1;B1=0;B0=1;S1=0;S0=1;
        #2 A3=1;A2=1;A1=0;A0=0;B3=1;B2=1;B1=1;B0=0;S1=0;S0=1;
        #2 A3=1;A2=1;A1=0;A0=0;B3=1;B2=1;B1=1;B0=1;S1=0;S0=1;
        #2 A3=1;A2=1;A1=0;A0=1;B3=0;B2=0;B1=0;B0=0;S1=0;S0=1;
        #2 A3=1;A2=1;A1=0;A0=1;B3=0;B2=0;B1=0;B0=1;S1=0;S0=1;
        #2 A3=1;A2=1;A1=0;A0=1;B3=0;B2=0;B1=1;B0=0;S1=0;S0=1;
        #2 A3=1;A2=1;A1=0;A0=1;B3=0;B2=0;B1=1;B0=1;S1=0;S0=1;
        #2 A3=1;A2=1;A1=0;A0=1;B3=0;B2=1;B1=0;B0=0;S1=0;S0=1;
        #2 A3=1;A2=1;A1=0;A0=1;B3=0;B2=1;B1=0;B0=1;S1=0;S0=1;
        #2 A3=1;A2=1;A1=0;A0=1;B3=0;B2=1;B1=1;B0=0;S1=0;S0=1;
        #2 A3=1;A2=1;A1=0;A0=1;B3=0;B2=1;B1=1;B0=1;S1=0;S0=1;
        #2 A3=1;A2=1;A1=0;A0=1;B3=1;B2=0;B1=0;B0=0;S1=0;S0=1;
        #2 A3=1;A2=1;A1=0;A0=1;B3=1;B2=0;B1=0;B0=1;S1=0;S0=1;
        #2 A3=1;A2=1;A1=0;A0=1;B3=1;B2=0;B1=1;B0=0;S1=0;S0=1;
        #2 A3=1;A2=1;A1=0;A0=1;B3=1;B2=0;B1=1;B0=1;S1=0;S0=1;
        #2 A3=1;A2=1;A1=0;A0=1;B3=1;B2=1;B1=0;B0=0;S1=0;S0=1;
        #2 A3=1;A2=1;A1=0;A0=1;B3=1;B2=1;B1=0;B0=1;S1=0;S0=1;
        #2 A3=1;A2=1;A1=0;A0=1;B3=1;B2=1;B1=1;B0=0;S1=0;S0=1;
        #2 A3=1;A2=1;A1=0;A0=1;B3=1;B2=1;B1=1;B0=1;S1=0;S0=1;
        #2 A3=1;A2=1;A1=1;A0=0;B3=0;B2=0;B1=0;B0=0;S1=0;S0=1;
        #2 A3=1;A2=1;A1=1;A0=0;B3=0;B2=0;B1=0;B0=1;S1=0;S0=1;
        #2 A3=1;A2=1;A1=1;A0=0;B3=0;B2=0;B1=1;B0=0;S1=0;S0=1;
        #2 A3=1;A2=1;A1=1;A0=0;B3=0;B2=0;B1=1;B0=1;S1=0;S0=1;
        #2 A3=1;A2=1;A1=1;A0=0;B3=0;B2=1;B1=0;B0=0;S1=0;S0=1;
        #2 A3=1;A2=1;A1=1;A0=0;B3=0;B2=1;B1=0;B0=1;S1=0;S0=1;
        #2 A3=1;A2=1;A1=1;A0=0;B3=0;B2=1;B1=1;B0=0;S1=0;S0=1;
        #2 A3=1;A2=1;A1=1;A0=0;B3=0;B2=1;B1=1;B0=1;S1=0;S0=1;
        #2 A3=1;A2=1;A1=1;A0=0;B3=1;B2=0;B1=0;B0=0;S1=0;S0=1;
        #2 A3=1;A2=1;A1=1;A0=0;B3=1;B2=0;B1=0;B0=1;S1=0;S0=1;
        #2 A3=1;A2=1;A1=1;A0=0;B3=1;B2=0;B1=1;B0=0;S1=0;S0=1;
        #2 A3=1;A2=1;A1=1;A0=0;B3=1;B2=0;B1=1;B0=1;S1=0;S0=1;
        #2 A3=1;A2=1;A1=1;A0=0;B3=1;B2=1;B1=0;B0=0;S1=0;S0=1;
        #2 A3=1;A2=1;A1=1;A0=0;B3=1;B2=1;B1=0;B0=1;S1=0;S0=1;
        #2 A3=1;A2=1;A1=1;A0=0;B3=1;B2=1;B1=1;B0=0;S1=0;S0=1;
        #2 A3=1;A2=1;A1=1;A0=0;B3=1;B2=1;B1=1;B0=1;S1=0;S0=1;
        #2 A3=1;A2=1;A1=1;A0=1;B3=0;B2=0;B1=0;B0=0;S1=0;S0=1;
        #2 A3=1;A2=1;A1=1;A0=1;B3=0;B2=0;B1=0;B0=1;S1=0;S0=1;
        #2 A3=1;A2=1;A1=1;A0=1;B3=0;B2=0;B1=1;B0=0;S1=0;S0=1;
        #2 A3=1;A2=1;A1=1;A0=1;B3=0;B2=0;B1=1;B0=1;S1=0;S0=1;
        #2 A3=1;A2=1;A1=1;A0=1;B3=0;B2=1;B1=0;B0=0;S1=0;S0=1;
        #2 A3=1;A2=1;A1=1;A0=1;B3=0;B2=1;B1=0;B0=1;S1=0;S0=1;
        #2 A3=1;A2=1;A1=1;A0=1;B3=0;B2=1;B1=1;B0=0;S1=0;S0=1;
        #2 A3=1;A2=1;A1=1;A0=1;B3=0;B2=1;B1=1;B0=1;S1=0;S0=1;
        #2 A3=1;A2=1;A1=1;A0=1;B3=1;B2=0;B1=0;B0=0;S1=0;S0=1;
        #2 A3=1;A2=1;A1=1;A0=1;B3=1;B2=0;B1=0;B0=1;S1=0;S0=1;
        #2 A3=1;A2=1;A1=1;A0=1;B3=1;B2=0;B1=1;B0=0;S1=0;S0=1;
        #2 A3=1;A2=1;A1=1;A0=1;B3=1;B2=0;B1=1;B0=1;S1=0;S0=1;
        #2 A3=1;A2=1;A1=1;A0=1;B3=1;B2=1;B1=0;B0=0;S1=0;S0=1;
        #2 A3=1;A2=1;A1=1;A0=1;B3=1;B2=1;B1=0;B0=1;S1=0;S0=1;
        #2 A3=1;A2=1;A1=1;A0=1;B3=1;B2=1;B1=1;B0=0;S1=0;S0=1;
        #2 A3=1;A2=1;A1=1;A0=1;B3=1;B2=1;B1=1;B0=1;S1=0;S0=1;
        #2 A3=0;A2=0;A1=0;A0=0;B3=0;B2=0;B1=0;B0=0;S1=1;S0=0;
        #2 A3=0;A2=0;A1=0;A0=0;B3=0;B2=0;B1=0;B0=1;S1=1;S0=0;
        #2 A3=0;A2=0;A1=0;A0=0;B3=0;B2=0;B1=1;B0=0;S1=1;S0=0;
        #2 A3=0;A2=0;A1=0;A0=0;B3=0;B2=0;B1=1;B0=1;S1=1;S0=0;
        #2 A3=0;A2=0;A1=0;A0=0;B3=0;B2=1;B1=0;B0=0;S1=1;S0=0;
        #2 A3=0;A2=0;A1=0;A0=0;B3=0;B2=1;B1=0;B0=1;S1=1;S0=0;
        #2 A3=0;A2=0;A1=0;A0=0;B3=0;B2=1;B1=1;B0=0;S1=1;S0=0;
        #2 A3=0;A2=0;A1=0;A0=0;B3=0;B2=1;B1=1;B0=1;S1=1;S0=0;
        #2 A3=0;A2=0;A1=0;A0=0;B3=1;B2=0;B1=0;B0=0;S1=1;S0=0;
        #2 A3=0;A2=0;A1=0;A0=0;B3=1;B2=0;B1=0;B0=1;S1=1;S0=0;
        #2 A3=0;A2=0;A1=0;A0=0;B3=1;B2=0;B1=1;B0=0;S1=1;S0=0;
        #2 A3=0;A2=0;A1=0;A0=0;B3=1;B2=0;B1=1;B0=1;S1=1;S0=0;
        #2 A3=0;A2=0;A1=0;A0=0;B3=1;B2=1;B1=0;B0=0;S1=1;S0=0;
        #2 A3=0;A2=0;A1=0;A0=0;B3=1;B2=1;B1=0;B0=1;S1=1;S0=0;
        #2 A3=0;A2=0;A1=0;A0=0;B3=1;B2=1;B1=1;B0=0;S1=1;S0=0;
        #2 A3=0;A2=0;A1=0;A0=0;B3=1;B2=1;B1=1;B0=1;S1=1;S0=0;
        #2 A3=0;A2=0;A1=0;A0=1;B3=0;B2=0;B1=0;B0=0;S1=1;S0=0;
        #2 A3=0;A2=0;A1=0;A0=1;B3=0;B2=0;B1=0;B0=1;S1=1;S0=0;
        #2 A3=0;A2=0;A1=0;A0=1;B3=0;B2=0;B1=1;B0=0;S1=1;S0=0;
        #2 A3=0;A2=0;A1=0;A0=1;B3=0;B2=0;B1=1;B0=1;S1=1;S0=0;
        #2 A3=0;A2=0;A1=0;A0=1;B3=0;B2=1;B1=0;B0=0;S1=1;S0=0;
        #2 A3=0;A2=0;A1=0;A0=1;B3=0;B2=1;B1=0;B0=1;S1=1;S0=0;
        #2 A3=0;A2=0;A1=0;A0=1;B3=0;B2=1;B1=1;B0=0;S1=1;S0=0;
        #2 A3=0;A2=0;A1=0;A0=1;B3=0;B2=1;B1=1;B0=1;S1=1;S0=0;
        #2 A3=0;A2=0;A1=0;A0=1;B3=1;B2=0;B1=0;B0=0;S1=1;S0=0;
        #2 A3=0;A2=0;A1=0;A0=1;B3=1;B2=0;B1=0;B0=1;S1=1;S0=0;
        #2 A3=0;A2=0;A1=0;A0=1;B3=1;B2=0;B1=1;B0=0;S1=1;S0=0;
        #2 A3=0;A2=0;A1=0;A0=1;B3=1;B2=0;B1=1;B0=1;S1=1;S0=0;
        #2 A3=0;A2=0;A1=0;A0=1;B3=1;B2=1;B1=0;B0=0;S1=1;S0=0;
        #2 A3=0;A2=0;A1=0;A0=1;B3=1;B2=1;B1=0;B0=1;S1=1;S0=0;
        #2 A3=0;A2=0;A1=0;A0=1;B3=1;B2=1;B1=1;B0=0;S1=1;S0=0;
        #2 A3=0;A2=0;A1=0;A0=1;B3=1;B2=1;B1=1;B0=1;S1=1;S0=0;
        #2 A3=0;A2=0;A1=1;A0=0;B3=0;B2=0;B1=0;B0=0;S1=1;S0=0;
        #2 A3=0;A2=0;A1=1;A0=0;B3=0;B2=0;B1=0;B0=1;S1=1;S0=0;
        #2 A3=0;A2=0;A1=1;A0=0;B3=0;B2=0;B1=1;B0=0;S1=1;S0=0;
        #2 A3=0;A2=0;A1=1;A0=0;B3=0;B2=0;B1=1;B0=1;S1=1;S0=0;
        #2 A3=0;A2=0;A1=1;A0=0;B3=0;B2=1;B1=0;B0=0;S1=1;S0=0;
        #2 A3=0;A2=0;A1=1;A0=0;B3=0;B2=1;B1=0;B0=1;S1=1;S0=0;
        #2 A3=0;A2=0;A1=1;A0=0;B3=0;B2=1;B1=1;B0=0;S1=1;S0=0;
        #2 A3=0;A2=0;A1=1;A0=0;B3=0;B2=1;B1=1;B0=1;S1=1;S0=0;
        #2 A3=0;A2=0;A1=1;A0=0;B3=1;B2=0;B1=0;B0=0;S1=1;S0=0;
        #2 A3=0;A2=0;A1=1;A0=0;B3=1;B2=0;B1=0;B0=1;S1=1;S0=0;
        #2 A3=0;A2=0;A1=1;A0=0;B3=1;B2=0;B1=1;B0=0;S1=1;S0=0;
        #2 A3=0;A2=0;A1=1;A0=0;B3=1;B2=0;B1=1;B0=1;S1=1;S0=0;
        #2 A3=0;A2=0;A1=1;A0=0;B3=1;B2=1;B1=0;B0=0;S1=1;S0=0;
        #2 A3=0;A2=0;A1=1;A0=0;B3=1;B2=1;B1=0;B0=1;S1=1;S0=0;
        #2 A3=0;A2=0;A1=1;A0=0;B3=1;B2=1;B1=1;B0=0;S1=1;S0=0;
        #2 A3=0;A2=0;A1=1;A0=0;B3=1;B2=1;B1=1;B0=1;S1=1;S0=0;
        #2 A3=0;A2=0;A1=1;A0=1;B3=0;B2=0;B1=0;B0=0;S1=1;S0=0;
        #2 A3=0;A2=0;A1=1;A0=1;B3=0;B2=0;B1=0;B0=1;S1=1;S0=0;
        #2 A3=0;A2=0;A1=1;A0=1;B3=0;B2=0;B1=1;B0=0;S1=1;S0=0;
        #2 A3=0;A2=0;A1=1;A0=1;B3=0;B2=0;B1=1;B0=1;S1=1;S0=0;
        #2 A3=0;A2=0;A1=1;A0=1;B3=0;B2=1;B1=0;B0=0;S1=1;S0=0;
        #2 A3=0;A2=0;A1=1;A0=1;B3=0;B2=1;B1=0;B0=1;S1=1;S0=0;
        #2 A3=0;A2=0;A1=1;A0=1;B3=0;B2=1;B1=1;B0=0;S1=1;S0=0;
        #2 A3=0;A2=0;A1=1;A0=1;B3=0;B2=1;B1=1;B0=1;S1=1;S0=0;
        #2 A3=0;A2=0;A1=1;A0=1;B3=1;B2=0;B1=0;B0=0;S1=1;S0=0;
        #2 A3=0;A2=0;A1=1;A0=1;B3=1;B2=0;B1=0;B0=1;S1=1;S0=0;
        #2 A3=0;A2=0;A1=1;A0=1;B3=1;B2=0;B1=1;B0=0;S1=1;S0=0;
        #2 A3=0;A2=0;A1=1;A0=1;B3=1;B2=0;B1=1;B0=1;S1=1;S0=0;
        #2 A3=0;A2=0;A1=1;A0=1;B3=1;B2=1;B1=0;B0=0;S1=1;S0=0;
        #2 A3=0;A2=0;A1=1;A0=1;B3=1;B2=1;B1=0;B0=1;S1=1;S0=0;
        #2 A3=0;A2=0;A1=1;A0=1;B3=1;B2=1;B1=1;B0=0;S1=1;S0=0;
        #2 A3=0;A2=0;A1=1;A0=1;B3=1;B2=1;B1=1;B0=1;S1=1;S0=0;
        #2 A3=0;A2=1;A1=0;A0=0;B3=0;B2=0;B1=0;B0=0;S1=1;S0=0;
        #2 A3=0;A2=1;A1=0;A0=0;B3=0;B2=0;B1=0;B0=1;S1=1;S0=0;
        #2 A3=0;A2=1;A1=0;A0=0;B3=0;B2=0;B1=1;B0=0;S1=1;S0=0;
        #2 A3=0;A2=1;A1=0;A0=0;B3=0;B2=0;B1=1;B0=1;S1=1;S0=0;
        #2 A3=0;A2=1;A1=0;A0=0;B3=0;B2=1;B1=0;B0=0;S1=1;S0=0;
        #2 A3=0;A2=1;A1=0;A0=0;B3=0;B2=1;B1=0;B0=1;S1=1;S0=0;
        #2 A3=0;A2=1;A1=0;A0=0;B3=0;B2=1;B1=1;B0=0;S1=1;S0=0;
        #2 A3=0;A2=1;A1=0;A0=0;B3=0;B2=1;B1=1;B0=1;S1=1;S0=0;
        #2 A3=0;A2=1;A1=0;A0=0;B3=1;B2=0;B1=0;B0=0;S1=1;S0=0;
        #2 A3=0;A2=1;A1=0;A0=0;B3=1;B2=0;B1=0;B0=1;S1=1;S0=0;
        #2 A3=0;A2=1;A1=0;A0=0;B3=1;B2=0;B1=1;B0=0;S1=1;S0=0;
        #2 A3=0;A2=1;A1=0;A0=0;B3=1;B2=0;B1=1;B0=1;S1=1;S0=0;
        #2 A3=0;A2=1;A1=0;A0=0;B3=1;B2=1;B1=0;B0=0;S1=1;S0=0;
        #2 A3=0;A2=1;A1=0;A0=0;B3=1;B2=1;B1=0;B0=1;S1=1;S0=0;
        #2 A3=0;A2=1;A1=0;A0=0;B3=1;B2=1;B1=1;B0=0;S1=1;S0=0;
        #2 A3=0;A2=1;A1=0;A0=0;B3=1;B2=1;B1=1;B0=1;S1=1;S0=0;
        #2 A3=0;A2=1;A1=0;A0=1;B3=0;B2=0;B1=0;B0=0;S1=1;S0=0;
        #2 A3=0;A2=1;A1=0;A0=1;B3=0;B2=0;B1=0;B0=1;S1=1;S0=0;
        #2 A3=0;A2=1;A1=0;A0=1;B3=0;B2=0;B1=1;B0=0;S1=1;S0=0;
        #2 A3=0;A2=1;A1=0;A0=1;B3=0;B2=0;B1=1;B0=1;S1=1;S0=0;
        #2 A3=0;A2=1;A1=0;A0=1;B3=0;B2=1;B1=0;B0=0;S1=1;S0=0;
        #2 A3=0;A2=1;A1=0;A0=1;B3=0;B2=1;B1=0;B0=1;S1=1;S0=0;
        #2 A3=0;A2=1;A1=0;A0=1;B3=0;B2=1;B1=1;B0=0;S1=1;S0=0;
        #2 A3=0;A2=1;A1=0;A0=1;B3=0;B2=1;B1=1;B0=1;S1=1;S0=0;
        #2 A3=0;A2=1;A1=0;A0=1;B3=1;B2=0;B1=0;B0=0;S1=1;S0=0;
        #2 A3=0;A2=1;A1=0;A0=1;B3=1;B2=0;B1=0;B0=1;S1=1;S0=0;
        #2 A3=0;A2=1;A1=0;A0=1;B3=1;B2=0;B1=1;B0=0;S1=1;S0=0;
        #2 A3=0;A2=1;A1=0;A0=1;B3=1;B2=0;B1=1;B0=1;S1=1;S0=0;
        #2 A3=0;A2=1;A1=0;A0=1;B3=1;B2=1;B1=0;B0=0;S1=1;S0=0;
        #2 A3=0;A2=1;A1=0;A0=1;B3=1;B2=1;B1=0;B0=1;S1=1;S0=0;
        #2 A3=0;A2=1;A1=0;A0=1;B3=1;B2=1;B1=1;B0=0;S1=1;S0=0;
        #2 A3=0;A2=1;A1=0;A0=1;B3=1;B2=1;B1=1;B0=1;S1=1;S0=0;
        #2 A3=0;A2=1;A1=1;A0=0;B3=0;B2=0;B1=0;B0=0;S1=1;S0=0;
        #2 A3=0;A2=1;A1=1;A0=0;B3=0;B2=0;B1=0;B0=1;S1=1;S0=0;
        #2 A3=0;A2=1;A1=1;A0=0;B3=0;B2=0;B1=1;B0=0;S1=1;S0=0;
        #2 A3=0;A2=1;A1=1;A0=0;B3=0;B2=0;B1=1;B0=1;S1=1;S0=0;
        #2 A3=0;A2=1;A1=1;A0=0;B3=0;B2=1;B1=0;B0=0;S1=1;S0=0;
        #2 A3=0;A2=1;A1=1;A0=0;B3=0;B2=1;B1=0;B0=1;S1=1;S0=0;
        #2 A3=0;A2=1;A1=1;A0=0;B3=0;B2=1;B1=1;B0=0;S1=1;S0=0;
        #2 A3=0;A2=1;A1=1;A0=0;B3=0;B2=1;B1=1;B0=1;S1=1;S0=0;
        #2 A3=0;A2=1;A1=1;A0=0;B3=1;B2=0;B1=0;B0=0;S1=1;S0=0;
        #2 A3=0;A2=1;A1=1;A0=0;B3=1;B2=0;B1=0;B0=1;S1=1;S0=0;
        #2 A3=0;A2=1;A1=1;A0=0;B3=1;B2=0;B1=1;B0=0;S1=1;S0=0;
        #2 A3=0;A2=1;A1=1;A0=0;B3=1;B2=0;B1=1;B0=1;S1=1;S0=0;
        #2 A3=0;A2=1;A1=1;A0=0;B3=1;B2=1;B1=0;B0=0;S1=1;S0=0;
        #2 A3=0;A2=1;A1=1;A0=0;B3=1;B2=1;B1=0;B0=1;S1=1;S0=0;
        #2 A3=0;A2=1;A1=1;A0=0;B3=1;B2=1;B1=1;B0=0;S1=1;S0=0;
        #2 A3=0;A2=1;A1=1;A0=0;B3=1;B2=1;B1=1;B0=1;S1=1;S0=0;
        #2 A3=0;A2=1;A1=1;A0=1;B3=0;B2=0;B1=0;B0=0;S1=1;S0=0;
        #2 A3=0;A2=1;A1=1;A0=1;B3=0;B2=0;B1=0;B0=1;S1=1;S0=0;
        #2 A3=0;A2=1;A1=1;A0=1;B3=0;B2=0;B1=1;B0=0;S1=1;S0=0;
        #2 A3=0;A2=1;A1=1;A0=1;B3=0;B2=0;B1=1;B0=1;S1=1;S0=0;
        #2 A3=0;A2=1;A1=1;A0=1;B3=0;B2=1;B1=0;B0=0;S1=1;S0=0;
        #2 A3=0;A2=1;A1=1;A0=1;B3=0;B2=1;B1=0;B0=1;S1=1;S0=0;
        #2 A3=0;A2=1;A1=1;A0=1;B3=0;B2=1;B1=1;B0=0;S1=1;S0=0;
        #2 A3=0;A2=1;A1=1;A0=1;B3=0;B2=1;B1=1;B0=1;S1=1;S0=0;
        #2 A3=0;A2=1;A1=1;A0=1;B3=1;B2=0;B1=0;B0=0;S1=1;S0=0;
        #2 A3=0;A2=1;A1=1;A0=1;B3=1;B2=0;B1=0;B0=1;S1=1;S0=0;
        #2 A3=0;A2=1;A1=1;A0=1;B3=1;B2=0;B1=1;B0=0;S1=1;S0=0;
        #2 A3=0;A2=1;A1=1;A0=1;B3=1;B2=0;B1=1;B0=1;S1=1;S0=0;
        #2 A3=0;A2=1;A1=1;A0=1;B3=1;B2=1;B1=0;B0=0;S1=1;S0=0;
        #2 A3=0;A2=1;A1=1;A0=1;B3=1;B2=1;B1=0;B0=1;S1=1;S0=0;
        #2 A3=0;A2=1;A1=1;A0=1;B3=1;B2=1;B1=1;B0=0;S1=1;S0=0;
        #2 A3=0;A2=1;A1=1;A0=1;B3=1;B2=1;B1=1;B0=1;S1=1;S0=0;
        #2 A3=1;A2=0;A1=0;A0=0;B3=0;B2=0;B1=0;B0=0;S1=1;S0=0;
        #2 A3=1;A2=0;A1=0;A0=0;B3=0;B2=0;B1=0;B0=1;S1=1;S0=0;
        #2 A3=1;A2=0;A1=0;A0=0;B3=0;B2=0;B1=1;B0=0;S1=1;S0=0;
        #2 A3=1;A2=0;A1=0;A0=0;B3=0;B2=0;B1=1;B0=1;S1=1;S0=0;
        #2 A3=1;A2=0;A1=0;A0=0;B3=0;B2=1;B1=0;B0=0;S1=1;S0=0;
        #2 A3=1;A2=0;A1=0;A0=0;B3=0;B2=1;B1=0;B0=1;S1=1;S0=0;
        #2 A3=1;A2=0;A1=0;A0=0;B3=0;B2=1;B1=1;B0=0;S1=1;S0=0;
        #2 A3=1;A2=0;A1=0;A0=0;B3=0;B2=1;B1=1;B0=1;S1=1;S0=0;
        #2 A3=1;A2=0;A1=0;A0=0;B3=1;B2=0;B1=0;B0=0;S1=1;S0=0;
        #2 A3=1;A2=0;A1=0;A0=0;B3=1;B2=0;B1=0;B0=1;S1=1;S0=0;
        #2 A3=1;A2=0;A1=0;A0=0;B3=1;B2=0;B1=1;B0=0;S1=1;S0=0;
        #2 A3=1;A2=0;A1=0;A0=0;B3=1;B2=0;B1=1;B0=1;S1=1;S0=0;
        #2 A3=1;A2=0;A1=0;A0=0;B3=1;B2=1;B1=0;B0=0;S1=1;S0=0;
        #2 A3=1;A2=0;A1=0;A0=0;B3=1;B2=1;B1=0;B0=1;S1=1;S0=0;
        #2 A3=1;A2=0;A1=0;A0=0;B3=1;B2=1;B1=1;B0=0;S1=1;S0=0;
        #2 A3=1;A2=0;A1=0;A0=0;B3=1;B2=1;B1=1;B0=1;S1=1;S0=0;
        #2 A3=1;A2=0;A1=0;A0=1;B3=0;B2=0;B1=0;B0=0;S1=1;S0=0;
        #2 A3=1;A2=0;A1=0;A0=1;B3=0;B2=0;B1=0;B0=1;S1=1;S0=0;
        #2 A3=1;A2=0;A1=0;A0=1;B3=0;B2=0;B1=1;B0=0;S1=1;S0=0;
        #2 A3=1;A2=0;A1=0;A0=1;B3=0;B2=0;B1=1;B0=1;S1=1;S0=0;
        #2 A3=1;A2=0;A1=0;A0=1;B3=0;B2=1;B1=0;B0=0;S1=1;S0=0;
        #2 A3=1;A2=0;A1=0;A0=1;B3=0;B2=1;B1=0;B0=1;S1=1;S0=0;
        #2 A3=1;A2=0;A1=0;A0=1;B3=0;B2=1;B1=1;B0=0;S1=1;S0=0;
        #2 A3=1;A2=0;A1=0;A0=1;B3=0;B2=1;B1=1;B0=1;S1=1;S0=0;
        #2 A3=1;A2=0;A1=0;A0=1;B3=1;B2=0;B1=0;B0=0;S1=1;S0=0;
        #2 A3=1;A2=0;A1=0;A0=1;B3=1;B2=0;B1=0;B0=1;S1=1;S0=0;
        #2 A3=1;A2=0;A1=0;A0=1;B3=1;B2=0;B1=1;B0=0;S1=1;S0=0;
        #2 A3=1;A2=0;A1=0;A0=1;B3=1;B2=0;B1=1;B0=1;S1=1;S0=0;
        #2 A3=1;A2=0;A1=0;A0=1;B3=1;B2=1;B1=0;B0=0;S1=1;S0=0;
        #2 A3=1;A2=0;A1=0;A0=1;B3=1;B2=1;B1=0;B0=1;S1=1;S0=0;
        #2 A3=1;A2=0;A1=0;A0=1;B3=1;B2=1;B1=1;B0=0;S1=1;S0=0;
        #2 A3=1;A2=0;A1=0;A0=1;B3=1;B2=1;B1=1;B0=1;S1=1;S0=0;
        #2 A3=1;A2=0;A1=1;A0=0;B3=0;B2=0;B1=0;B0=0;S1=1;S0=0;
        #2 A3=1;A2=0;A1=1;A0=0;B3=0;B2=0;B1=0;B0=1;S1=1;S0=0;
        #2 A3=1;A2=0;A1=1;A0=0;B3=0;B2=0;B1=1;B0=0;S1=1;S0=0;
        #2 A3=1;A2=0;A1=1;A0=0;B3=0;B2=0;B1=1;B0=1;S1=1;S0=0;
        #2 A3=1;A2=0;A1=1;A0=0;B3=0;B2=1;B1=0;B0=0;S1=1;S0=0;
        #2 A3=1;A2=0;A1=1;A0=0;B3=0;B2=1;B1=0;B0=1;S1=1;S0=0;
        #2 A3=1;A2=0;A1=1;A0=0;B3=0;B2=1;B1=1;B0=0;S1=1;S0=0;
        #2 A3=1;A2=0;A1=1;A0=0;B3=0;B2=1;B1=1;B0=1;S1=1;S0=0;
        #2 A3=1;A2=0;A1=1;A0=0;B3=1;B2=0;B1=0;B0=0;S1=1;S0=0;
        #2 A3=1;A2=0;A1=1;A0=0;B3=1;B2=0;B1=0;B0=1;S1=1;S0=0;
        #2 A3=1;A2=0;A1=1;A0=0;B3=1;B2=0;B1=1;B0=0;S1=1;S0=0;
        #2 A3=1;A2=0;A1=1;A0=0;B3=1;B2=0;B1=1;B0=1;S1=1;S0=0;
        #2 A3=1;A2=0;A1=1;A0=0;B3=1;B2=1;B1=0;B0=0;S1=1;S0=0;
        #2 A3=1;A2=0;A1=1;A0=0;B3=1;B2=1;B1=0;B0=1;S1=1;S0=0;
        #2 A3=1;A2=0;A1=1;A0=0;B3=1;B2=1;B1=1;B0=0;S1=1;S0=0;
        #2 A3=1;A2=0;A1=1;A0=0;B3=1;B2=1;B1=1;B0=1;S1=1;S0=0;
        #2 A3=1;A2=0;A1=1;A0=1;B3=0;B2=0;B1=0;B0=0;S1=1;S0=0;
        #2 A3=1;A2=0;A1=1;A0=1;B3=0;B2=0;B1=0;B0=1;S1=1;S0=0;
        #2 A3=1;A2=0;A1=1;A0=1;B3=0;B2=0;B1=1;B0=0;S1=1;S0=0;
        #2 A3=1;A2=0;A1=1;A0=1;B3=0;B2=0;B1=1;B0=1;S1=1;S0=0;
        #2 A3=1;A2=0;A1=1;A0=1;B3=0;B2=1;B1=0;B0=0;S1=1;S0=0;
        #2 A3=1;A2=0;A1=1;A0=1;B3=0;B2=1;B1=0;B0=1;S1=1;S0=0;
        #2 A3=1;A2=0;A1=1;A0=1;B3=0;B2=1;B1=1;B0=0;S1=1;S0=0;
        #2 A3=1;A2=0;A1=1;A0=1;B3=0;B2=1;B1=1;B0=1;S1=1;S0=0;
        #2 A3=1;A2=0;A1=1;A0=1;B3=1;B2=0;B1=0;B0=0;S1=1;S0=0;
        #2 A3=1;A2=0;A1=1;A0=1;B3=1;B2=0;B1=0;B0=1;S1=1;S0=0;
        #2 A3=1;A2=0;A1=1;A0=1;B3=1;B2=0;B1=1;B0=0;S1=1;S0=0;
        #2 A3=1;A2=0;A1=1;A0=1;B3=1;B2=0;B1=1;B0=1;S1=1;S0=0;
        #2 A3=1;A2=0;A1=1;A0=1;B3=1;B2=1;B1=0;B0=0;S1=1;S0=0;
        #2 A3=1;A2=0;A1=1;A0=1;B3=1;B2=1;B1=0;B0=1;S1=1;S0=0;
        #2 A3=1;A2=0;A1=1;A0=1;B3=1;B2=1;B1=1;B0=0;S1=1;S0=0;
        #2 A3=1;A2=0;A1=1;A0=1;B3=1;B2=1;B1=1;B0=1;S1=1;S0=0;
        #2 A3=1;A2=1;A1=0;A0=0;B3=0;B2=0;B1=0;B0=0;S1=1;S0=0;
        #2 A3=1;A2=1;A1=0;A0=0;B3=0;B2=0;B1=0;B0=1;S1=1;S0=0;
        #2 A3=1;A2=1;A1=0;A0=0;B3=0;B2=0;B1=1;B0=0;S1=1;S0=0;
        #2 A3=1;A2=1;A1=0;A0=0;B3=0;B2=0;B1=1;B0=1;S1=1;S0=0;
        #2 A3=1;A2=1;A1=0;A0=0;B3=0;B2=1;B1=0;B0=0;S1=1;S0=0;
        #2 A3=1;A2=1;A1=0;A0=0;B3=0;B2=1;B1=0;B0=1;S1=1;S0=0;
        #2 A3=1;A2=1;A1=0;A0=0;B3=0;B2=1;B1=1;B0=0;S1=1;S0=0;
        #2 A3=1;A2=1;A1=0;A0=0;B3=0;B2=1;B1=1;B0=1;S1=1;S0=0;
        #2 A3=1;A2=1;A1=0;A0=0;B3=1;B2=0;B1=0;B0=0;S1=1;S0=0;
        #2 A3=1;A2=1;A1=0;A0=0;B3=1;B2=0;B1=0;B0=1;S1=1;S0=0;
        #2 A3=1;A2=1;A1=0;A0=0;B3=1;B2=0;B1=1;B0=0;S1=1;S0=0;
        #2 A3=1;A2=1;A1=0;A0=0;B3=1;B2=0;B1=1;B0=1;S1=1;S0=0;
        #2 A3=1;A2=1;A1=0;A0=0;B3=1;B2=1;B1=0;B0=0;S1=1;S0=0;
        #2 A3=1;A2=1;A1=0;A0=0;B3=1;B2=1;B1=0;B0=1;S1=1;S0=0;
        #2 A3=1;A2=1;A1=0;A0=0;B3=1;B2=1;B1=1;B0=0;S1=1;S0=0;
        #2 A3=1;A2=1;A1=0;A0=0;B3=1;B2=1;B1=1;B0=1;S1=1;S0=0;
        #2 A3=1;A2=1;A1=0;A0=1;B3=0;B2=0;B1=0;B0=0;S1=1;S0=0;
        #2 A3=1;A2=1;A1=0;A0=1;B3=0;B2=0;B1=0;B0=1;S1=1;S0=0;
        #2 A3=1;A2=1;A1=0;A0=1;B3=0;B2=0;B1=1;B0=0;S1=1;S0=0;
        #2 A3=1;A2=1;A1=0;A0=1;B3=0;B2=0;B1=1;B0=1;S1=1;S0=0;
        #2 A3=1;A2=1;A1=0;A0=1;B3=0;B2=1;B1=0;B0=0;S1=1;S0=0;
        #2 A3=1;A2=1;A1=0;A0=1;B3=0;B2=1;B1=0;B0=1;S1=1;S0=0;
        #2 A3=1;A2=1;A1=0;A0=1;B3=0;B2=1;B1=1;B0=0;S1=1;S0=0;
        #2 A3=1;A2=1;A1=0;A0=1;B3=0;B2=1;B1=1;B0=1;S1=1;S0=0;
        #2 A3=1;A2=1;A1=0;A0=1;B3=1;B2=0;B1=0;B0=0;S1=1;S0=0;
        #2 A3=1;A2=1;A1=0;A0=1;B3=1;B2=0;B1=0;B0=1;S1=1;S0=0;
        #2 A3=1;A2=1;A1=0;A0=1;B3=1;B2=0;B1=1;B0=0;S1=1;S0=0;
        #2 A3=1;A2=1;A1=0;A0=1;B3=1;B2=0;B1=1;B0=1;S1=1;S0=0;
        #2 A3=1;A2=1;A1=0;A0=1;B3=1;B2=1;B1=0;B0=0;S1=1;S0=0;
        #2 A3=1;A2=1;A1=0;A0=1;B3=1;B2=1;B1=0;B0=1;S1=1;S0=0;
        #2 A3=1;A2=1;A1=0;A0=1;B3=1;B2=1;B1=1;B0=0;S1=1;S0=0;
        #2 A3=1;A2=1;A1=0;A0=1;B3=1;B2=1;B1=1;B0=1;S1=1;S0=0;
        #2 A3=1;A2=1;A1=1;A0=0;B3=0;B2=0;B1=0;B0=0;S1=1;S0=0;
        #2 A3=1;A2=1;A1=1;A0=0;B3=0;B2=0;B1=0;B0=1;S1=1;S0=0;
        #2 A3=1;A2=1;A1=1;A0=0;B3=0;B2=0;B1=1;B0=0;S1=1;S0=0;
        #2 A3=1;A2=1;A1=1;A0=0;B3=0;B2=0;B1=1;B0=1;S1=1;S0=0;
        #2 A3=1;A2=1;A1=1;A0=0;B3=0;B2=1;B1=0;B0=0;S1=1;S0=0;
        #2 A3=1;A2=1;A1=1;A0=0;B3=0;B2=1;B1=0;B0=1;S1=1;S0=0;
        #2 A3=1;A2=1;A1=1;A0=0;B3=0;B2=1;B1=1;B0=0;S1=1;S0=0;
        #2 A3=1;A2=1;A1=1;A0=0;B3=0;B2=1;B1=1;B0=1;S1=1;S0=0;
        #2 A3=1;A2=1;A1=1;A0=0;B3=1;B2=0;B1=0;B0=0;S1=1;S0=0;
        #2 A3=1;A2=1;A1=1;A0=0;B3=1;B2=0;B1=0;B0=1;S1=1;S0=0;
        #2 A3=1;A2=1;A1=1;A0=0;B3=1;B2=0;B1=1;B0=0;S1=1;S0=0;
        #2 A3=1;A2=1;A1=1;A0=0;B3=1;B2=0;B1=1;B0=1;S1=1;S0=0;
        #2 A3=1;A2=1;A1=1;A0=0;B3=1;B2=1;B1=0;B0=0;S1=1;S0=0;
        #2 A3=1;A2=1;A1=1;A0=0;B3=1;B2=1;B1=0;B0=1;S1=1;S0=0;
        #2 A3=1;A2=1;A1=1;A0=0;B3=1;B2=1;B1=1;B0=0;S1=1;S0=0;
        #2 A3=1;A2=1;A1=1;A0=0;B3=1;B2=1;B1=1;B0=1;S1=1;S0=0;
        #2 A3=1;A2=1;A1=1;A0=1;B3=0;B2=0;B1=0;B0=0;S1=1;S0=0;
        #2 A3=1;A2=1;A1=1;A0=1;B3=0;B2=0;B1=0;B0=1;S1=1;S0=0;
        #2 A3=1;A2=1;A1=1;A0=1;B3=0;B2=0;B1=1;B0=0;S1=1;S0=0;
        #2 A3=1;A2=1;A1=1;A0=1;B3=0;B2=0;B1=1;B0=1;S1=1;S0=0;
        #2 A3=1;A2=1;A1=1;A0=1;B3=0;B2=1;B1=0;B0=0;S1=1;S0=0;
        #2 A3=1;A2=1;A1=1;A0=1;B3=0;B2=1;B1=0;B0=1;S1=1;S0=0;
        #2 A3=1;A2=1;A1=1;A0=1;B3=0;B2=1;B1=1;B0=0;S1=1;S0=0;
        #2 A3=1;A2=1;A1=1;A0=1;B3=0;B2=1;B1=1;B0=1;S1=1;S0=0;
        #2 A3=1;A2=1;A1=1;A0=1;B3=1;B2=0;B1=0;B0=0;S1=1;S0=0;
        #2 A3=1;A2=1;A1=1;A0=1;B3=1;B2=0;B1=0;B0=1;S1=1;S0=0;
        #2 A3=1;A2=1;A1=1;A0=1;B3=1;B2=0;B1=1;B0=0;S1=1;S0=0;
        #2 A3=1;A2=1;A1=1;A0=1;B3=1;B2=0;B1=1;B0=1;S1=1;S0=0;
        #2 A3=1;A2=1;A1=1;A0=1;B3=1;B2=1;B1=0;B0=0;S1=1;S0=0;
        #2 A3=1;A2=1;A1=1;A0=1;B3=1;B2=1;B1=0;B0=1;S1=1;S0=0;
        #2 A3=1;A2=1;A1=1;A0=1;B3=1;B2=1;B1=1;B0=0;S1=1;S0=0;
        #2 A3=1;A2=1;A1=1;A0=1;B3=1;B2=1;B1=1;B0=1;S1=1;S0=0;
        #2 A3=0;A2=0;A1=0;A0=0;B3=0;B2=0;B1=0;B0=0;S1=1;S0=1;
        #2 A3=0;A2=0;A1=0;A0=0;B3=0;B2=0;B1=0;B0=1;S1=1;S0=1;
        #2 A3=0;A2=0;A1=0;A0=0;B3=0;B2=0;B1=1;B0=0;S1=1;S0=1;
        #2 A3=0;A2=0;A1=0;A0=0;B3=0;B2=0;B1=1;B0=1;S1=1;S0=1;
        #2 A3=0;A2=0;A1=0;A0=0;B3=0;B2=1;B1=0;B0=0;S1=1;S0=1;
        #2 A3=0;A2=0;A1=0;A0=0;B3=0;B2=1;B1=0;B0=1;S1=1;S0=1;
        #2 A3=0;A2=0;A1=0;A0=0;B3=0;B2=1;B1=1;B0=0;S1=1;S0=1;
        #2 A3=0;A2=0;A1=0;A0=0;B3=0;B2=1;B1=1;B0=1;S1=1;S0=1;
        #2 A3=0;A2=0;A1=0;A0=0;B3=1;B2=0;B1=0;B0=0;S1=1;S0=1;
        #2 A3=0;A2=0;A1=0;A0=0;B3=1;B2=0;B1=0;B0=1;S1=1;S0=1;
        #2 A3=0;A2=0;A1=0;A0=0;B3=1;B2=0;B1=1;B0=0;S1=1;S0=1;
        #2 A3=0;A2=0;A1=0;A0=0;B3=1;B2=0;B1=1;B0=1;S1=1;S0=1;
        #2 A3=0;A2=0;A1=0;A0=0;B3=1;B2=1;B1=0;B0=0;S1=1;S0=1;
        #2 A3=0;A2=0;A1=0;A0=0;B3=1;B2=1;B1=0;B0=1;S1=1;S0=1;
        #2 A3=0;A2=0;A1=0;A0=0;B3=1;B2=1;B1=1;B0=0;S1=1;S0=1;
        #2 A3=0;A2=0;A1=0;A0=0;B3=1;B2=1;B1=1;B0=1;S1=1;S0=1;
        #2 A3=0;A2=0;A1=0;A0=1;B3=0;B2=0;B1=0;B0=0;S1=1;S0=1;
        #2 A3=0;A2=0;A1=0;A0=1;B3=0;B2=0;B1=0;B0=1;S1=1;S0=1;
        #2 A3=0;A2=0;A1=0;A0=1;B3=0;B2=0;B1=1;B0=0;S1=1;S0=1;
        #2 A3=0;A2=0;A1=0;A0=1;B3=0;B2=0;B1=1;B0=1;S1=1;S0=1;
        #2 A3=0;A2=0;A1=0;A0=1;B3=0;B2=1;B1=0;B0=0;S1=1;S0=1;
        #2 A3=0;A2=0;A1=0;A0=1;B3=0;B2=1;B1=0;B0=1;S1=1;S0=1;
        #2 A3=0;A2=0;A1=0;A0=1;B3=0;B2=1;B1=1;B0=0;S1=1;S0=1;
        #2 A3=0;A2=0;A1=0;A0=1;B3=0;B2=1;B1=1;B0=1;S1=1;S0=1;
        #2 A3=0;A2=0;A1=0;A0=1;B3=1;B2=0;B1=0;B0=0;S1=1;S0=1;
        #2 A3=0;A2=0;A1=0;A0=1;B3=1;B2=0;B1=0;B0=1;S1=1;S0=1;
        #2 A3=0;A2=0;A1=0;A0=1;B3=1;B2=0;B1=1;B0=0;S1=1;S0=1;
        #2 A3=0;A2=0;A1=0;A0=1;B3=1;B2=0;B1=1;B0=1;S1=1;S0=1;
        #2 A3=0;A2=0;A1=0;A0=1;B3=1;B2=1;B1=0;B0=0;S1=1;S0=1;
        #2 A3=0;A2=0;A1=0;A0=1;B3=1;B2=1;B1=0;B0=1;S1=1;S0=1;
        #2 A3=0;A2=0;A1=0;A0=1;B3=1;B2=1;B1=1;B0=0;S1=1;S0=1;
        #2 A3=0;A2=0;A1=0;A0=1;B3=1;B2=1;B1=1;B0=1;S1=1;S0=1;
        #2 A3=0;A2=0;A1=1;A0=0;B3=0;B2=0;B1=0;B0=0;S1=1;S0=1;
        #2 A3=0;A2=0;A1=1;A0=0;B3=0;B2=0;B1=0;B0=1;S1=1;S0=1;
        #2 A3=0;A2=0;A1=1;A0=0;B3=0;B2=0;B1=1;B0=0;S1=1;S0=1;
        #2 A3=0;A2=0;A1=1;A0=0;B3=0;B2=0;B1=1;B0=1;S1=1;S0=1;
        #2 A3=0;A2=0;A1=1;A0=0;B3=0;B2=1;B1=0;B0=0;S1=1;S0=1;
        #2 A3=0;A2=0;A1=1;A0=0;B3=0;B2=1;B1=0;B0=1;S1=1;S0=1;
        #2 A3=0;A2=0;A1=1;A0=0;B3=0;B2=1;B1=1;B0=0;S1=1;S0=1;
        #2 A3=0;A2=0;A1=1;A0=0;B3=0;B2=1;B1=1;B0=1;S1=1;S0=1;
        #2 A3=0;A2=0;A1=1;A0=0;B3=1;B2=0;B1=0;B0=0;S1=1;S0=1;
        #2 A3=0;A2=0;A1=1;A0=0;B3=1;B2=0;B1=0;B0=1;S1=1;S0=1;
        #2 A3=0;A2=0;A1=1;A0=0;B3=1;B2=0;B1=1;B0=0;S1=1;S0=1;
        #2 A3=0;A2=0;A1=1;A0=0;B3=1;B2=0;B1=1;B0=1;S1=1;S0=1;
        #2 A3=0;A2=0;A1=1;A0=0;B3=1;B2=1;B1=0;B0=0;S1=1;S0=1;
        #2 A3=0;A2=0;A1=1;A0=0;B3=1;B2=1;B1=0;B0=1;S1=1;S0=1;
        #2 A3=0;A2=0;A1=1;A0=0;B3=1;B2=1;B1=1;B0=0;S1=1;S0=1;
        #2 A3=0;A2=0;A1=1;A0=0;B3=1;B2=1;B1=1;B0=1;S1=1;S0=1;
        #2 A3=0;A2=0;A1=1;A0=1;B3=0;B2=0;B1=0;B0=0;S1=1;S0=1;
        #2 A3=0;A2=0;A1=1;A0=1;B3=0;B2=0;B1=0;B0=1;S1=1;S0=1;
        #2 A3=0;A2=0;A1=1;A0=1;B3=0;B2=0;B1=1;B0=0;S1=1;S0=1;
        #2 A3=0;A2=0;A1=1;A0=1;B3=0;B2=0;B1=1;B0=1;S1=1;S0=1;
        #2 A3=0;A2=0;A1=1;A0=1;B3=0;B2=1;B1=0;B0=0;S1=1;S0=1;
        #2 A3=0;A2=0;A1=1;A0=1;B3=0;B2=1;B1=0;B0=1;S1=1;S0=1;
        #2 A3=0;A2=0;A1=1;A0=1;B3=0;B2=1;B1=1;B0=0;S1=1;S0=1;
        #2 A3=0;A2=0;A1=1;A0=1;B3=0;B2=1;B1=1;B0=1;S1=1;S0=1;
        #2 A3=0;A2=0;A1=1;A0=1;B3=1;B2=0;B1=0;B0=0;S1=1;S0=1;
        #2 A3=0;A2=0;A1=1;A0=1;B3=1;B2=0;B1=0;B0=1;S1=1;S0=1;
        #2 A3=0;A2=0;A1=1;A0=1;B3=1;B2=0;B1=1;B0=0;S1=1;S0=1;
        #2 A3=0;A2=0;A1=1;A0=1;B3=1;B2=0;B1=1;B0=1;S1=1;S0=1;
        #2 A3=0;A2=0;A1=1;A0=1;B3=1;B2=1;B1=0;B0=0;S1=1;S0=1;
        #2 A3=0;A2=0;A1=1;A0=1;B3=1;B2=1;B1=0;B0=1;S1=1;S0=1;
        #2 A3=0;A2=0;A1=1;A0=1;B3=1;B2=1;B1=1;B0=0;S1=1;S0=1;
        #2 A3=0;A2=0;A1=1;A0=1;B3=1;B2=1;B1=1;B0=1;S1=1;S0=1;
        #2 A3=0;A2=1;A1=0;A0=0;B3=0;B2=0;B1=0;B0=0;S1=1;S0=1;
        #2 A3=0;A2=1;A1=0;A0=0;B3=0;B2=0;B1=0;B0=1;S1=1;S0=1;
        #2 A3=0;A2=1;A1=0;A0=0;B3=0;B2=0;B1=1;B0=0;S1=1;S0=1;
        #2 A3=0;A2=1;A1=0;A0=0;B3=0;B2=0;B1=1;B0=1;S1=1;S0=1;
        #2 A3=0;A2=1;A1=0;A0=0;B3=0;B2=1;B1=0;B0=0;S1=1;S0=1;
        #2 A3=0;A2=1;A1=0;A0=0;B3=0;B2=1;B1=0;B0=1;S1=1;S0=1;
        #2 A3=0;A2=1;A1=0;A0=0;B3=0;B2=1;B1=1;B0=0;S1=1;S0=1;
        #2 A3=0;A2=1;A1=0;A0=0;B3=0;B2=1;B1=1;B0=1;S1=1;S0=1;
        #2 A3=0;A2=1;A1=0;A0=0;B3=1;B2=0;B1=0;B0=0;S1=1;S0=1;
        #2 A3=0;A2=1;A1=0;A0=0;B3=1;B2=0;B1=0;B0=1;S1=1;S0=1;
        #2 A3=0;A2=1;A1=0;A0=0;B3=1;B2=0;B1=1;B0=0;S1=1;S0=1;
        #2 A3=0;A2=1;A1=0;A0=0;B3=1;B2=0;B1=1;B0=1;S1=1;S0=1;
        #2 A3=0;A2=1;A1=0;A0=0;B3=1;B2=1;B1=0;B0=0;S1=1;S0=1;
        #2 A3=0;A2=1;A1=0;A0=0;B3=1;B2=1;B1=0;B0=1;S1=1;S0=1;
        #2 A3=0;A2=1;A1=0;A0=0;B3=1;B2=1;B1=1;B0=0;S1=1;S0=1;
        #2 A3=0;A2=1;A1=0;A0=0;B3=1;B2=1;B1=1;B0=1;S1=1;S0=1;
        #2 A3=0;A2=1;A1=0;A0=1;B3=0;B2=0;B1=0;B0=0;S1=1;S0=1;
        #2 A3=0;A2=1;A1=0;A0=1;B3=0;B2=0;B1=0;B0=1;S1=1;S0=1;
        #2 A3=0;A2=1;A1=0;A0=1;B3=0;B2=0;B1=1;B0=0;S1=1;S0=1;
        #2 A3=0;A2=1;A1=0;A0=1;B3=0;B2=0;B1=1;B0=1;S1=1;S0=1;
        #2 A3=0;A2=1;A1=0;A0=1;B3=0;B2=1;B1=0;B0=0;S1=1;S0=1;
        #2 A3=0;A2=1;A1=0;A0=1;B3=0;B2=1;B1=0;B0=1;S1=1;S0=1;
        #2 A3=0;A2=1;A1=0;A0=1;B3=0;B2=1;B1=1;B0=0;S1=1;S0=1;
        #2 A3=0;A2=1;A1=0;A0=1;B3=0;B2=1;B1=1;B0=1;S1=1;S0=1;
        #2 A3=0;A2=1;A1=0;A0=1;B3=1;B2=0;B1=0;B0=0;S1=1;S0=1;
        #2 A3=0;A2=1;A1=0;A0=1;B3=1;B2=0;B1=0;B0=1;S1=1;S0=1;
        #2 A3=0;A2=1;A1=0;A0=1;B3=1;B2=0;B1=1;B0=0;S1=1;S0=1;
        #2 A3=0;A2=1;A1=0;A0=1;B3=1;B2=0;B1=1;B0=1;S1=1;S0=1;
        #2 A3=0;A2=1;A1=0;A0=1;B3=1;B2=1;B1=0;B0=0;S1=1;S0=1;
        #2 A3=0;A2=1;A1=0;A0=1;B3=1;B2=1;B1=0;B0=1;S1=1;S0=1;
        #2 A3=0;A2=1;A1=0;A0=1;B3=1;B2=1;B1=1;B0=0;S1=1;S0=1;
        #2 A3=0;A2=1;A1=0;A0=1;B3=1;B2=1;B1=1;B0=1;S1=1;S0=1;
        #2 A3=0;A2=1;A1=1;A0=0;B3=0;B2=0;B1=0;B0=0;S1=1;S0=1;
        #2 A3=0;A2=1;A1=1;A0=0;B3=0;B2=0;B1=0;B0=1;S1=1;S0=1;
        #2 A3=0;A2=1;A1=1;A0=0;B3=0;B2=0;B1=1;B0=0;S1=1;S0=1;
        #2 A3=0;A2=1;A1=1;A0=0;B3=0;B2=0;B1=1;B0=1;S1=1;S0=1;
        #2 A3=0;A2=1;A1=1;A0=0;B3=0;B2=1;B1=0;B0=0;S1=1;S0=1;
        #2 A3=0;A2=1;A1=1;A0=0;B3=0;B2=1;B1=0;B0=1;S1=1;S0=1;
        #2 A3=0;A2=1;A1=1;A0=0;B3=0;B2=1;B1=1;B0=0;S1=1;S0=1;
        #2 A3=0;A2=1;A1=1;A0=0;B3=0;B2=1;B1=1;B0=1;S1=1;S0=1;
        #2 A3=0;A2=1;A1=1;A0=0;B3=1;B2=0;B1=0;B0=0;S1=1;S0=1;
        #2 A3=0;A2=1;A1=1;A0=0;B3=1;B2=0;B1=0;B0=1;S1=1;S0=1;
        #2 A3=0;A2=1;A1=1;A0=0;B3=1;B2=0;B1=1;B0=0;S1=1;S0=1;
        #2 A3=0;A2=1;A1=1;A0=0;B3=1;B2=0;B1=1;B0=1;S1=1;S0=1;
        #2 A3=0;A2=1;A1=1;A0=0;B3=1;B2=1;B1=0;B0=0;S1=1;S0=1;
        #2 A3=0;A2=1;A1=1;A0=0;B3=1;B2=1;B1=0;B0=1;S1=1;S0=1;
        #2 A3=0;A2=1;A1=1;A0=0;B3=1;B2=1;B1=1;B0=0;S1=1;S0=1;
        #2 A3=0;A2=1;A1=1;A0=0;B3=1;B2=1;B1=1;B0=1;S1=1;S0=1;
        #2 A3=0;A2=1;A1=1;A0=1;B3=0;B2=0;B1=0;B0=0;S1=1;S0=1;
        #2 A3=0;A2=1;A1=1;A0=1;B3=0;B2=0;B1=0;B0=1;S1=1;S0=1;
        #2 A3=0;A2=1;A1=1;A0=1;B3=0;B2=0;B1=1;B0=0;S1=1;S0=1;
        #2 A3=0;A2=1;A1=1;A0=1;B3=0;B2=0;B1=1;B0=1;S1=1;S0=1;
        #2 A3=0;A2=1;A1=1;A0=1;B3=0;B2=1;B1=0;B0=0;S1=1;S0=1;
        #2 A3=0;A2=1;A1=1;A0=1;B3=0;B2=1;B1=0;B0=1;S1=1;S0=1;
        #2 A3=0;A2=1;A1=1;A0=1;B3=0;B2=1;B1=1;B0=0;S1=1;S0=1;
        #2 A3=0;A2=1;A1=1;A0=1;B3=0;B2=1;B1=1;B0=1;S1=1;S0=1;
        #2 A3=0;A2=1;A1=1;A0=1;B3=1;B2=0;B1=0;B0=0;S1=1;S0=1;
        #2 A3=0;A2=1;A1=1;A0=1;B3=1;B2=0;B1=0;B0=1;S1=1;S0=1;
        #2 A3=0;A2=1;A1=1;A0=1;B3=1;B2=0;B1=1;B0=0;S1=1;S0=1;
        #2 A3=0;A2=1;A1=1;A0=1;B3=1;B2=0;B1=1;B0=1;S1=1;S0=1;
        #2 A3=0;A2=1;A1=1;A0=1;B3=1;B2=1;B1=0;B0=0;S1=1;S0=1;
        #2 A3=0;A2=1;A1=1;A0=1;B3=1;B2=1;B1=0;B0=1;S1=1;S0=1;
        #2 A3=0;A2=1;A1=1;A0=1;B3=1;B2=1;B1=1;B0=0;S1=1;S0=1;
        #2 A3=0;A2=1;A1=1;A0=1;B3=1;B2=1;B1=1;B0=1;S1=1;S0=1;
        #2 A3=1;A2=0;A1=0;A0=0;B3=0;B2=0;B1=0;B0=0;S1=1;S0=1;
        #2 A3=1;A2=0;A1=0;A0=0;B3=0;B2=0;B1=0;B0=1;S1=1;S0=1;
        #2 A3=1;A2=0;A1=0;A0=0;B3=0;B2=0;B1=1;B0=0;S1=1;S0=1;
        #2 A3=1;A2=0;A1=0;A0=0;B3=0;B2=0;B1=1;B0=1;S1=1;S0=1;
        #2 A3=1;A2=0;A1=0;A0=0;B3=0;B2=1;B1=0;B0=0;S1=1;S0=1;
        #2 A3=1;A2=0;A1=0;A0=0;B3=0;B2=1;B1=0;B0=1;S1=1;S0=1;
        #2 A3=1;A2=0;A1=0;A0=0;B3=0;B2=1;B1=1;B0=0;S1=1;S0=1;
        #2 A3=1;A2=0;A1=0;A0=0;B3=0;B2=1;B1=1;B0=1;S1=1;S0=1;
        #2 A3=1;A2=0;A1=0;A0=0;B3=1;B2=0;B1=0;B0=0;S1=1;S0=1;
        #2 A3=1;A2=0;A1=0;A0=0;B3=1;B2=0;B1=0;B0=1;S1=1;S0=1;
        #2 A3=1;A2=0;A1=0;A0=0;B3=1;B2=0;B1=1;B0=0;S1=1;S0=1;
        #2 A3=1;A2=0;A1=0;A0=0;B3=1;B2=0;B1=1;B0=1;S1=1;S0=1;
        #2 A3=1;A2=0;A1=0;A0=0;B3=1;B2=1;B1=0;B0=0;S1=1;S0=1;
        #2 A3=1;A2=0;A1=0;A0=0;B3=1;B2=1;B1=0;B0=1;S1=1;S0=1;
        #2 A3=1;A2=0;A1=0;A0=0;B3=1;B2=1;B1=1;B0=0;S1=1;S0=1;
        #2 A3=1;A2=0;A1=0;A0=0;B3=1;B2=1;B1=1;B0=1;S1=1;S0=1;
        #2 A3=1;A2=0;A1=0;A0=1;B3=0;B2=0;B1=0;B0=0;S1=1;S0=1;
        #2 A3=1;A2=0;A1=0;A0=1;B3=0;B2=0;B1=0;B0=1;S1=1;S0=1;
        #2 A3=1;A2=0;A1=0;A0=1;B3=0;B2=0;B1=1;B0=0;S1=1;S0=1;
        #2 A3=1;A2=0;A1=0;A0=1;B3=0;B2=0;B1=1;B0=1;S1=1;S0=1;
        #2 A3=1;A2=0;A1=0;A0=1;B3=0;B2=1;B1=0;B0=0;S1=1;S0=1;
        #2 A3=1;A2=0;A1=0;A0=1;B3=0;B2=1;B1=0;B0=1;S1=1;S0=1;
        #2 A3=1;A2=0;A1=0;A0=1;B3=0;B2=1;B1=1;B0=0;S1=1;S0=1;
        #2 A3=1;A2=0;A1=0;A0=1;B3=0;B2=1;B1=1;B0=1;S1=1;S0=1;
        #2 A3=1;A2=0;A1=0;A0=1;B3=1;B2=0;B1=0;B0=0;S1=1;S0=1;
        #2 A3=1;A2=0;A1=0;A0=1;B3=1;B2=0;B1=0;B0=1;S1=1;S0=1;
        #2 A3=1;A2=0;A1=0;A0=1;B3=1;B2=0;B1=1;B0=0;S1=1;S0=1;
        #2 A3=1;A2=0;A1=0;A0=1;B3=1;B2=0;B1=1;B0=1;S1=1;S0=1;
        #2 A3=1;A2=0;A1=0;A0=1;B3=1;B2=1;B1=0;B0=0;S1=1;S0=1;
        #2 A3=1;A2=0;A1=0;A0=1;B3=1;B2=1;B1=0;B0=1;S1=1;S0=1;
        #2 A3=1;A2=0;A1=0;A0=1;B3=1;B2=1;B1=1;B0=0;S1=1;S0=1;
        #2 A3=1;A2=0;A1=0;A0=1;B3=1;B2=1;B1=1;B0=1;S1=1;S0=1;
        #2 A3=1;A2=0;A1=1;A0=0;B3=0;B2=0;B1=0;B0=0;S1=1;S0=1;
        #2 A3=1;A2=0;A1=1;A0=0;B3=0;B2=0;B1=0;B0=1;S1=1;S0=1;
        #2 A3=1;A2=0;A1=1;A0=0;B3=0;B2=0;B1=1;B0=0;S1=1;S0=1;
        #2 A3=1;A2=0;A1=1;A0=0;B3=0;B2=0;B1=1;B0=1;S1=1;S0=1;
        #2 A3=1;A2=0;A1=1;A0=0;B3=0;B2=1;B1=0;B0=0;S1=1;S0=1;
        #2 A3=1;A2=0;A1=1;A0=0;B3=0;B2=1;B1=0;B0=1;S1=1;S0=1;
        #2 A3=1;A2=0;A1=1;A0=0;B3=0;B2=1;B1=1;B0=0;S1=1;S0=1;
        #2 A3=1;A2=0;A1=1;A0=0;B3=0;B2=1;B1=1;B0=1;S1=1;S0=1;
        #2 A3=1;A2=0;A1=1;A0=0;B3=1;B2=0;B1=0;B0=0;S1=1;S0=1;
        #2 A3=1;A2=0;A1=1;A0=0;B3=1;B2=0;B1=0;B0=1;S1=1;S0=1;
        #2 A3=1;A2=0;A1=1;A0=0;B3=1;B2=0;B1=1;B0=0;S1=1;S0=1;
        #2 A3=1;A2=0;A1=1;A0=0;B3=1;B2=0;B1=1;B0=1;S1=1;S0=1;
        #2 A3=1;A2=0;A1=1;A0=0;B3=1;B2=1;B1=0;B0=0;S1=1;S0=1;
        #2 A3=1;A2=0;A1=1;A0=0;B3=1;B2=1;B1=0;B0=1;S1=1;S0=1;
        #2 A3=1;A2=0;A1=1;A0=0;B3=1;B2=1;B1=1;B0=0;S1=1;S0=1;
        #2 A3=1;A2=0;A1=1;A0=0;B3=1;B2=1;B1=1;B0=1;S1=1;S0=1;
        #2 A3=1;A2=0;A1=1;A0=1;B3=0;B2=0;B1=0;B0=0;S1=1;S0=1;
        #2 A3=1;A2=0;A1=1;A0=1;B3=0;B2=0;B1=0;B0=1;S1=1;S0=1;
        #2 A3=1;A2=0;A1=1;A0=1;B3=0;B2=0;B1=1;B0=0;S1=1;S0=1;
        #2 A3=1;A2=0;A1=1;A0=1;B3=0;B2=0;B1=1;B0=1;S1=1;S0=1;
        #2 A3=1;A2=0;A1=1;A0=1;B3=0;B2=1;B1=0;B0=0;S1=1;S0=1;
        #2 A3=1;A2=0;A1=1;A0=1;B3=0;B2=1;B1=0;B0=1;S1=1;S0=1;
        #2 A3=1;A2=0;A1=1;A0=1;B3=0;B2=1;B1=1;B0=0;S1=1;S0=1;
        #2 A3=1;A2=0;A1=1;A0=1;B3=0;B2=1;B1=1;B0=1;S1=1;S0=1;
        #2 A3=1;A2=0;A1=1;A0=1;B3=1;B2=0;B1=0;B0=0;S1=1;S0=1;
        #2 A3=1;A2=0;A1=1;A0=1;B3=1;B2=0;B1=0;B0=1;S1=1;S0=1;
        #2 A3=1;A2=0;A1=1;A0=1;B3=1;B2=0;B1=1;B0=0;S1=1;S0=1;
        #2 A3=1;A2=0;A1=1;A0=1;B3=1;B2=0;B1=1;B0=1;S1=1;S0=1;
        #2 A3=1;A2=0;A1=1;A0=1;B3=1;B2=1;B1=0;B0=0;S1=1;S0=1;
        #2 A3=1;A2=0;A1=1;A0=1;B3=1;B2=1;B1=0;B0=1;S1=1;S0=1;
        #2 A3=1;A2=0;A1=1;A0=1;B3=1;B2=1;B1=1;B0=0;S1=1;S0=1;
        #2 A3=1;A2=0;A1=1;A0=1;B3=1;B2=1;B1=1;B0=1;S1=1;S0=1;
        #2 A3=1;A2=1;A1=0;A0=0;B3=0;B2=0;B1=0;B0=0;S1=1;S0=1;
        #2 A3=1;A2=1;A1=0;A0=0;B3=0;B2=0;B1=0;B0=1;S1=1;S0=1;
        #2 A3=1;A2=1;A1=0;A0=0;B3=0;B2=0;B1=1;B0=0;S1=1;S0=1;
        #2 A3=1;A2=1;A1=0;A0=0;B3=0;B2=0;B1=1;B0=1;S1=1;S0=1;
        #2 A3=1;A2=1;A1=0;A0=0;B3=0;B2=1;B1=0;B0=0;S1=1;S0=1;
        #2 A3=1;A2=1;A1=0;A0=0;B3=0;B2=1;B1=0;B0=1;S1=1;S0=1;
        #2 A3=1;A2=1;A1=0;A0=0;B3=0;B2=1;B1=1;B0=0;S1=1;S0=1;
        #2 A3=1;A2=1;A1=0;A0=0;B3=0;B2=1;B1=1;B0=1;S1=1;S0=1;
        #2 A3=1;A2=1;A1=0;A0=0;B3=1;B2=0;B1=0;B0=0;S1=1;S0=1;
        #2 A3=1;A2=1;A1=0;A0=0;B3=1;B2=0;B1=0;B0=1;S1=1;S0=1;
        #2 A3=1;A2=1;A1=0;A0=0;B3=1;B2=0;B1=1;B0=0;S1=1;S0=1;
        #2 A3=1;A2=1;A1=0;A0=0;B3=1;B2=0;B1=1;B0=1;S1=1;S0=1;
        #2 A3=1;A2=1;A1=0;A0=0;B3=1;B2=1;B1=0;B0=0;S1=1;S0=1;
        #2 A3=1;A2=1;A1=0;A0=0;B3=1;B2=1;B1=0;B0=1;S1=1;S0=1;
        #2 A3=1;A2=1;A1=0;A0=0;B3=1;B2=1;B1=1;B0=0;S1=1;S0=1;
        #2 A3=1;A2=1;A1=0;A0=0;B3=1;B2=1;B1=1;B0=1;S1=1;S0=1;
        #2 A3=1;A2=1;A1=0;A0=1;B3=0;B2=0;B1=0;B0=0;S1=1;S0=1;
        #2 A3=1;A2=1;A1=0;A0=1;B3=0;B2=0;B1=0;B0=1;S1=1;S0=1;
        #2 A3=1;A2=1;A1=0;A0=1;B3=0;B2=0;B1=1;B0=0;S1=1;S0=1;
        #2 A3=1;A2=1;A1=0;A0=1;B3=0;B2=0;B1=1;B0=1;S1=1;S0=1;
        #2 A3=1;A2=1;A1=0;A0=1;B3=0;B2=1;B1=0;B0=0;S1=1;S0=1;
        #2 A3=1;A2=1;A1=0;A0=1;B3=0;B2=1;B1=0;B0=1;S1=1;S0=1;
        #2 A3=1;A2=1;A1=0;A0=1;B3=0;B2=1;B1=1;B0=0;S1=1;S0=1;
        #2 A3=1;A2=1;A1=0;A0=1;B3=0;B2=1;B1=1;B0=1;S1=1;S0=1;
        #2 A3=1;A2=1;A1=0;A0=1;B3=1;B2=0;B1=0;B0=0;S1=1;S0=1;
        #2 A3=1;A2=1;A1=0;A0=1;B3=1;B2=0;B1=0;B0=1;S1=1;S0=1;
        #2 A3=1;A2=1;A1=0;A0=1;B3=1;B2=0;B1=1;B0=0;S1=1;S0=1;
        #2 A3=1;A2=1;A1=0;A0=1;B3=1;B2=0;B1=1;B0=1;S1=1;S0=1;
        #2 A3=1;A2=1;A1=0;A0=1;B3=1;B2=1;B1=0;B0=0;S1=1;S0=1;
        #2 A3=1;A2=1;A1=0;A0=1;B3=1;B2=1;B1=0;B0=1;S1=1;S0=1;
        #2 A3=1;A2=1;A1=0;A0=1;B3=1;B2=1;B1=1;B0=0;S1=1;S0=1;
        #2 A3=1;A2=1;A1=0;A0=1;B3=1;B2=1;B1=1;B0=1;S1=1;S0=1;
        #2 A3=1;A2=1;A1=1;A0=0;B3=0;B2=0;B1=0;B0=0;S1=1;S0=1;
        #2 A3=1;A2=1;A1=1;A0=0;B3=0;B2=0;B1=0;B0=1;S1=1;S0=1;
        #2 A3=1;A2=1;A1=1;A0=0;B3=0;B2=0;B1=1;B0=0;S1=1;S0=1;
        #2 A3=1;A2=1;A1=1;A0=0;B3=0;B2=0;B1=1;B0=1;S1=1;S0=1;
        #2 A3=1;A2=1;A1=1;A0=0;B3=0;B2=1;B1=0;B0=0;S1=1;S0=1;
        #2 A3=1;A2=1;A1=1;A0=0;B3=0;B2=1;B1=0;B0=1;S1=1;S0=1;
        #2 A3=1;A2=1;A1=1;A0=0;B3=0;B2=1;B1=1;B0=0;S1=1;S0=1;
        #2 A3=1;A2=1;A1=1;A0=0;B3=0;B2=1;B1=1;B0=1;S1=1;S0=1;
        #2 A3=1;A2=1;A1=1;A0=0;B3=1;B2=0;B1=0;B0=0;S1=1;S0=1;
        #2 A3=1;A2=1;A1=1;A0=0;B3=1;B2=0;B1=0;B0=1;S1=1;S0=1;
        #2 A3=1;A2=1;A1=1;A0=0;B3=1;B2=0;B1=1;B0=0;S1=1;S0=1;
        #2 A3=1;A2=1;A1=1;A0=0;B3=1;B2=0;B1=1;B0=1;S1=1;S0=1;
        #2 A3=1;A2=1;A1=1;A0=0;B3=1;B2=1;B1=0;B0=0;S1=1;S0=1;
        #2 A3=1;A2=1;A1=1;A0=0;B3=1;B2=1;B1=0;B0=1;S1=1;S0=1;
        #2 A3=1;A2=1;A1=1;A0=0;B3=1;B2=1;B1=1;B0=0;S1=1;S0=1;
        #2 A3=1;A2=1;A1=1;A0=0;B3=1;B2=1;B1=1;B0=1;S1=1;S0=1;
        #2 A3=1;A2=1;A1=1;A0=1;B3=0;B2=0;B1=0;B0=0;S1=1;S0=1;
        #2 A3=1;A2=1;A1=1;A0=1;B3=0;B2=0;B1=0;B0=1;S1=1;S0=1;
        #2 A3=1;A2=1;A1=1;A0=1;B3=0;B2=0;B1=1;B0=0;S1=1;S0=1;
        #2 A3=1;A2=1;A1=1;A0=1;B3=0;B2=0;B1=1;B0=1;S1=1;S0=1;
        #2 A3=1;A2=1;A1=1;A0=1;B3=0;B2=1;B1=0;B0=0;S1=1;S0=1;
        #2 A3=1;A2=1;A1=1;A0=1;B3=0;B2=1;B1=0;B0=1;S1=1;S0=1;
        #2 A3=1;A2=1;A1=1;A0=1;B3=0;B2=1;B1=1;B0=0;S1=1;S0=1;
        #2 A3=1;A2=1;A1=1;A0=1;B3=0;B2=1;B1=1;B0=1;S1=1;S0=1;
        #2 A3=1;A2=1;A1=1;A0=1;B3=1;B2=0;B1=0;B0=0;S1=1;S0=1;
        #2 A3=1;A2=1;A1=1;A0=1;B3=1;B2=0;B1=0;B0=1;S1=1;S0=1;
        #2 A3=1;A2=1;A1=1;A0=1;B3=1;B2=0;B1=1;B0=0;S1=1;S0=1;
        #2 A3=1;A2=1;A1=1;A0=1;B3=1;B2=0;B1=1;B0=1;S1=1;S0=1;
        #2 A3=1;A2=1;A1=1;A0=1;B3=1;B2=1;B1=0;B0=0;S1=1;S0=1;
        #2 A3=1;A2=1;A1=1;A0=1;B3=1;B2=1;B1=0;B0=1;S1=1;S0=1;
        #2 A3=1;A2=1;A1=1;A0=1;B3=1;B2=1;B1=1;B0=0;S1=1;S0=1;
        #2 A3=1;A2=1;A1=1;A0=1;B3=1;B2=1;B1=1;B0=1;S1=1;S0=1;
         #2 $finish;
    end 
endmodule