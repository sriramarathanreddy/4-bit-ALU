magic
tech scmos
timestamp 1701521160
<< nwell >>
rect 392 97 428 129
rect 448 97 484 129
rect 503 88 539 120
rect 590 97 626 129
rect 646 97 682 129
rect 701 88 737 120
rect 788 97 824 129
rect 844 97 880 129
rect 899 88 935 120
rect 986 97 1022 129
rect 1042 97 1078 129
rect 1097 88 1133 120
<< ntransistor >>
rect 435 51 439 71
rect 519 58 523 78
rect 633 51 637 71
rect 717 58 721 78
rect 831 51 835 71
rect 915 58 919 78
rect 1029 51 1033 71
rect 1113 58 1117 78
rect 435 11 439 31
rect 633 11 637 31
rect 831 11 835 31
rect 1029 11 1033 31
<< ptransistor >>
rect 409 103 411 123
rect 465 103 467 123
rect 520 94 522 114
rect 607 103 609 123
rect 663 103 665 123
rect 718 94 720 114
rect 805 103 807 123
rect 861 103 863 123
rect 916 94 918 114
rect 1003 103 1005 123
rect 1059 103 1061 123
rect 1114 94 1116 114
<< ndiffusion >>
rect 434 51 435 71
rect 439 51 440 71
rect 518 58 519 78
rect 523 58 524 78
rect 632 51 633 71
rect 637 51 638 71
rect 716 58 717 78
rect 721 58 722 78
rect 830 51 831 71
rect 835 51 836 71
rect 914 58 915 78
rect 919 58 920 78
rect 1028 51 1029 71
rect 1033 51 1034 71
rect 1112 58 1113 78
rect 1117 58 1118 78
rect 434 11 435 31
rect 439 11 440 31
rect 632 11 633 31
rect 637 11 638 31
rect 830 11 831 31
rect 835 11 836 31
rect 1028 11 1029 31
rect 1033 11 1034 31
<< pdiffusion >>
rect 408 103 409 123
rect 411 103 412 123
rect 464 103 465 123
rect 467 103 468 123
rect 519 94 520 114
rect 522 94 523 114
rect 606 103 607 123
rect 609 103 610 123
rect 662 103 663 123
rect 665 103 666 123
rect 717 94 718 114
rect 720 94 721 114
rect 804 103 805 123
rect 807 103 808 123
rect 860 103 861 123
rect 863 103 864 123
rect 915 94 916 114
rect 918 94 919 114
rect 1002 103 1003 123
rect 1005 103 1006 123
rect 1058 103 1059 123
rect 1061 103 1062 123
rect 1113 94 1114 114
rect 1116 94 1117 114
<< ndcontact >>
rect 424 51 434 71
rect 440 51 450 71
rect 508 58 518 78
rect 524 58 534 78
rect 622 51 632 71
rect 638 51 648 71
rect 706 58 716 78
rect 722 58 732 78
rect 820 51 830 71
rect 836 51 846 71
rect 904 58 914 78
rect 920 58 930 78
rect 1018 51 1028 71
rect 1034 51 1044 71
rect 1102 58 1112 78
rect 1118 58 1128 78
rect 424 11 434 31
rect 440 11 450 31
rect 622 11 632 31
rect 638 11 648 31
rect 820 11 830 31
rect 836 11 846 31
rect 1018 11 1028 31
rect 1034 11 1044 31
<< pdcontact >>
rect 398 103 408 123
rect 412 103 422 123
rect 454 103 464 123
rect 468 103 478 123
rect 509 94 519 114
rect 523 94 533 114
rect 596 103 606 123
rect 610 103 620 123
rect 652 103 662 123
rect 666 103 676 123
rect 707 94 717 114
rect 721 94 731 114
rect 794 103 804 123
rect 808 103 818 123
rect 850 103 860 123
rect 864 103 874 123
rect 905 94 915 114
rect 919 94 929 114
rect 992 103 1002 123
rect 1006 103 1016 123
rect 1048 103 1058 123
rect 1062 103 1072 123
rect 1103 94 1113 114
rect 1117 94 1127 114
<< psubstratepcontact >>
rect 392 1 396 5
rect 480 1 484 5
rect 503 1 507 5
rect 535 1 539 5
rect 590 1 594 5
rect 678 1 682 5
rect 701 1 705 5
rect 733 1 737 5
rect 788 1 792 5
rect 876 1 880 5
rect 899 1 903 5
rect 931 1 935 5
rect 986 1 990 5
rect 1074 1 1078 5
rect 1097 1 1101 5
rect 1129 1 1133 5
<< nsubstratencontact >>
rect 392 129 396 133
rect 480 129 484 133
rect 503 129 507 133
rect 535 129 539 133
rect 590 129 594 133
rect 678 129 682 133
rect 701 129 705 133
rect 733 129 737 133
rect 788 129 792 133
rect 876 129 880 133
rect 899 129 903 133
rect 931 129 935 133
rect 986 129 990 133
rect 1074 129 1078 133
rect 1097 129 1101 133
rect 1129 129 1133 133
<< polysilicon >>
rect 409 123 411 126
rect 465 123 467 126
rect 607 123 609 126
rect 663 123 665 126
rect 805 123 807 126
rect 861 123 863 126
rect 1003 123 1005 126
rect 1059 123 1061 126
rect 520 114 522 117
rect 409 94 411 103
rect 465 94 467 103
rect 718 114 720 117
rect 607 94 609 103
rect 663 94 665 103
rect 916 114 918 117
rect 805 94 807 103
rect 861 94 863 103
rect 1114 114 1116 117
rect 1003 94 1005 103
rect 1059 94 1061 103
rect 396 90 411 94
rect 452 90 467 94
rect 424 74 439 78
rect 435 71 439 74
rect 435 48 439 51
rect 463 38 467 90
rect 520 85 522 94
rect 594 90 609 94
rect 650 90 665 94
rect 505 83 522 85
rect 505 81 523 83
rect 519 78 523 81
rect 622 74 637 78
rect 633 71 637 74
rect 519 55 523 58
rect 633 48 637 51
rect 661 38 665 90
rect 718 85 720 94
rect 792 90 807 94
rect 848 90 863 94
rect 703 83 720 85
rect 703 81 721 83
rect 717 78 721 81
rect 820 74 835 78
rect 831 71 835 74
rect 717 55 721 58
rect 831 48 835 51
rect 859 38 863 90
rect 916 85 918 94
rect 990 90 1005 94
rect 1046 90 1061 94
rect 901 83 918 85
rect 901 81 919 83
rect 915 78 919 81
rect 1018 74 1033 78
rect 1029 71 1033 74
rect 915 55 919 58
rect 1029 48 1033 51
rect 1057 38 1061 90
rect 1114 85 1116 94
rect 1099 83 1116 85
rect 1099 81 1117 83
rect 1113 78 1117 81
rect 1113 55 1117 58
rect 424 34 467 38
rect 622 34 665 38
rect 820 34 863 38
rect 1018 34 1061 38
rect 435 31 439 34
rect 633 31 637 34
rect 831 31 835 34
rect 1029 31 1033 34
rect 435 8 439 11
rect 633 8 637 11
rect 831 8 835 11
rect 1029 8 1033 11
<< polycontact >>
rect 392 90 396 94
rect 420 74 424 78
rect 590 90 594 94
rect 501 81 505 85
rect 618 74 622 78
rect 788 90 792 94
rect 699 81 703 85
rect 816 74 820 78
rect 986 90 990 94
rect 897 81 901 85
rect 1014 74 1018 78
rect 1095 81 1099 85
rect 420 34 424 38
rect 618 34 622 38
rect 816 34 820 38
rect 1014 34 1018 38
<< metal1 >>
rect 396 129 480 133
rect 484 129 503 133
rect 507 129 535 133
rect 539 129 590 133
rect 594 129 678 133
rect 682 129 701 133
rect 705 129 733 133
rect 737 129 788 133
rect 792 129 876 133
rect 880 129 899 133
rect 903 129 931 133
rect 935 129 986 133
rect 990 129 1074 133
rect 1078 129 1097 133
rect 1101 129 1129 133
rect 398 123 408 129
rect 454 123 464 129
rect 377 90 392 94
rect 377 78 381 90
rect 412 85 422 103
rect 468 85 478 103
rect 509 114 519 129
rect 596 123 606 129
rect 652 123 662 129
rect 524 85 533 94
rect 575 90 590 94
rect 392 81 501 85
rect 524 81 547 85
rect 377 74 420 78
rect 440 71 450 81
rect 524 78 533 81
rect 575 78 579 90
rect 610 85 620 103
rect 666 85 676 103
rect 707 114 717 129
rect 794 123 804 129
rect 850 123 860 129
rect 722 85 731 94
rect 773 90 788 94
rect 590 81 699 85
rect 722 81 745 85
rect 575 74 618 78
rect 638 71 648 81
rect 722 78 731 81
rect 773 78 777 90
rect 808 85 818 103
rect 864 85 874 103
rect 905 114 915 129
rect 992 123 1002 129
rect 1048 123 1058 129
rect 920 85 929 94
rect 971 90 986 94
rect 788 81 897 85
rect 920 81 943 85
rect 424 45 434 51
rect 424 41 450 45
rect 405 34 420 38
rect 440 31 450 41
rect 424 5 434 11
rect 508 5 518 58
rect 773 74 816 78
rect 836 71 846 81
rect 920 78 929 81
rect 971 78 975 90
rect 1006 85 1016 103
rect 1062 85 1072 103
rect 1103 114 1113 129
rect 1118 85 1127 94
rect 986 81 1095 85
rect 1118 81 1141 85
rect 622 45 632 51
rect 622 41 648 45
rect 603 34 618 38
rect 638 31 648 41
rect 622 5 632 11
rect 706 5 716 58
rect 971 74 1014 78
rect 1034 71 1044 81
rect 1118 78 1127 81
rect 820 45 830 51
rect 820 41 846 45
rect 801 34 816 38
rect 836 31 846 41
rect 820 5 830 11
rect 904 5 914 58
rect 1018 45 1028 51
rect 1018 41 1044 45
rect 999 34 1014 38
rect 1034 31 1044 41
rect 1018 5 1028 11
rect 1102 5 1112 58
rect 396 1 480 5
rect 484 1 503 5
rect 507 1 535 5
rect 539 1 590 5
rect 594 1 678 5
rect 682 1 701 5
rect 705 1 733 5
rect 737 1 788 5
rect 792 1 876 5
rect 880 1 899 5
rect 903 1 931 5
rect 935 1 986 5
rect 990 1 1074 5
rect 1078 1 1097 5
rect 1101 1 1129 5
<< labels >>
rlabel metal1 392 1 1133 5 1 Gnd
rlabel metal1 392 129 1133 133 5 VDD
rlabel metal1 377 90 396 94 1 ANA0
rlabel metal1 575 90 594 94 1 ANA1
rlabel metal1 773 90 792 94 1 ANA2
rlabel metal1 971 90 990 94 1 ANA3
rlabel metal1 405 34 424 38 1 ANB0
rlabel metal1 603 34 622 38 1 ANB1
rlabel metal1 801 34 820 38 1 ANB2
rlabel metal1 999 34 1018 38 1 ANB3
rlabel metal1 533 81 547 85 1 OUT_AND0
rlabel metal1 731 81 745 85 1 OUT_AND1
rlabel metal1 929 81 943 85 1 OUT_AND2
rlabel metal1 1127 81 1141 85 1 OUT_AND3
<< end >>
