magic
tech scmos
timestamp 1701498759
<< nwell >>
rect 277 175 313 207
rect 333 175 369 207
rect 389 175 425 207
rect 445 175 481 207
rect 497 166 533 198
<< ntransistor >>
rect 320 129 324 149
rect 320 89 324 109
rect 320 49 324 69
rect 513 136 517 156
rect 320 10 324 30
<< ptransistor >>
rect 294 181 296 201
rect 350 181 352 201
rect 406 181 408 201
rect 462 181 464 201
rect 514 172 516 192
<< ndiffusion >>
rect 319 129 320 149
rect 324 129 325 149
rect 319 89 320 109
rect 324 89 325 109
rect 319 49 320 69
rect 324 49 325 69
rect 512 136 513 156
rect 517 136 518 156
rect 319 10 320 30
rect 324 10 325 30
<< pdiffusion >>
rect 293 181 294 201
rect 296 181 297 201
rect 349 181 350 201
rect 352 181 353 201
rect 405 181 406 201
rect 408 181 409 201
rect 461 181 462 201
rect 464 181 465 201
rect 513 172 514 192
rect 516 172 517 192
<< ndcontact >>
rect 309 129 319 149
rect 325 129 335 149
rect 309 89 319 109
rect 325 89 335 109
rect 309 49 319 69
rect 325 49 335 69
rect 502 136 512 156
rect 518 136 528 156
rect 309 10 319 30
rect 325 10 335 30
<< pdcontact >>
rect 283 181 293 201
rect 297 181 307 201
rect 339 181 349 201
rect 353 181 363 201
rect 395 181 405 201
rect 409 181 419 201
rect 451 181 461 201
rect 465 181 475 201
rect 503 172 513 192
rect 517 172 527 192
<< psubstratepcontact >>
rect 277 1 281 5
rect 477 1 481 5
rect 498 1 502 5
rect 530 1 534 5
<< nsubstratencontact >>
rect 277 207 281 211
rect 476 207 480 211
rect 498 207 502 211
rect 530 207 534 211
<< polysilicon >>
rect 294 201 296 204
rect 350 201 352 204
rect 406 201 408 204
rect 462 201 464 204
rect 514 192 516 195
rect 294 172 296 181
rect 350 172 352 181
rect 406 172 408 181
rect 462 172 464 181
rect 281 168 296 172
rect 337 168 352 172
rect 393 168 408 172
rect 449 168 464 172
rect 309 152 324 156
rect 320 149 324 152
rect 320 126 324 129
rect 348 116 352 168
rect 320 112 352 116
rect 320 109 324 112
rect 320 86 324 89
rect 404 76 408 168
rect 320 72 408 76
rect 320 69 324 72
rect 320 46 324 49
rect 460 37 464 168
rect 514 163 516 172
rect 499 161 516 163
rect 499 159 517 161
rect 513 156 517 159
rect 513 133 517 136
rect 320 33 464 37
rect 320 30 324 33
rect 320 7 324 10
<< polycontact >>
rect 277 168 281 172
rect 305 152 309 156
rect 316 112 320 116
rect 316 72 320 76
rect 495 159 499 163
rect 316 33 320 37
<< metal1 >>
rect 281 207 476 211
rect 480 207 498 211
rect 502 207 530 211
rect 283 201 293 207
rect 339 201 349 207
rect 395 201 405 207
rect 451 201 461 207
rect 262 168 277 172
rect 262 156 266 168
rect 297 163 307 181
rect 353 163 363 181
rect 409 163 419 181
rect 465 163 475 181
rect 503 192 513 207
rect 518 163 527 172
rect 277 159 495 163
rect 518 159 541 163
rect 262 152 305 156
rect 325 149 335 159
rect 518 156 527 159
rect 309 123 319 129
rect 309 119 335 123
rect 301 112 316 116
rect 325 109 335 119
rect 309 83 319 89
rect 309 79 335 83
rect 301 72 316 76
rect 325 69 335 79
rect 309 44 319 49
rect 309 40 335 44
rect 301 33 316 37
rect 325 30 335 40
rect 309 5 319 10
rect 502 5 512 136
rect 281 1 477 5
rect 481 1 498 5
rect 502 1 530 5
<< labels >>
rlabel metal1 262 168 281 172 1 A
rlabel metal1 277 207 534 211 5 VDD
rlabel metal1 522 159 541 163 1 OUT
rlabel metal1 277 1 534 5 1 Gnd
rlabel metal1 301 112 320 116 1 B
rlabel metal1 301 72 320 76 1 C
rlabel metal1 301 33 320 37 1 D
<< end >>
