magic
tech scmos
timestamp 1701500029
<< nwell >>
rect 0 0 36 32
rect 56 0 92 32
<< ntransistor >>
rect 43 -46 47 -26
rect 43 -86 47 -66
<< ptransistor >>
rect 17 6 19 26
rect 73 6 75 26
<< ndiffusion >>
rect 42 -46 43 -26
rect 47 -46 48 -26
rect 42 -86 43 -66
rect 47 -86 48 -66
<< pdiffusion >>
rect 16 6 17 26
rect 19 6 20 26
rect 72 6 73 26
rect 75 6 76 26
<< ndcontact >>
rect 32 -46 42 -26
rect 48 -46 58 -26
rect 32 -86 42 -66
rect 48 -86 58 -66
<< pdcontact >>
rect 6 6 16 26
rect 20 6 30 26
rect 62 6 72 26
rect 76 6 86 26
<< psubstratepcontact >>
rect 0 -96 4 -92
rect 88 -96 92 -92
<< nsubstratencontact >>
rect 0 32 4 36
rect 88 32 92 36
<< polysilicon >>
rect 17 26 19 29
rect 73 26 75 29
rect 17 -3 19 6
rect 73 -3 75 6
rect 4 -7 19 -3
rect 60 -7 75 -3
rect 32 -23 47 -19
rect 43 -26 47 -23
rect 43 -49 47 -46
rect 71 -59 75 -7
rect 32 -63 75 -59
rect 43 -66 47 -63
rect 43 -89 47 -86
<< polycontact >>
rect 0 -7 4 -3
rect 28 -23 32 -19
rect 28 -63 32 -59
<< metal1 >>
rect 4 32 88 36
rect 6 26 16 32
rect 62 26 72 32
rect -15 -7 0 -3
rect -15 -19 -11 -7
rect 20 -12 30 6
rect 76 -12 86 6
rect 0 -16 92 -12
rect -15 -23 28 -19
rect 48 -26 58 -16
rect 32 -52 42 -46
rect 32 -56 58 -52
rect 13 -63 28 -59
rect 48 -66 58 -56
rect 32 -92 42 -86
rect 4 -96 88 -92
<< labels >>
rlabel metal1 0 -96 92 -92 1 Gnd
rlabel metal1 0 -16 92 -12 1 OUT
rlabel metal1 0 32 92 36 5 VDD
rlabel metal1 -15 -7 4 -3 1 A
rlabel metal1 13 -63 32 -59 1 B
<< end >>
