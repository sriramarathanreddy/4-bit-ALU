* SPICE3 file created from comparator.ext - technology: scmos

.include TSMC_180nm.txt
.param SUPPLY = 1.8
.global Gnd
Vdd VDD Gnd 'SUPPLY'
.option scale=0.09u

VinCOA3 COA3 Gnd DC 0
VinCOA2 COA2 Gnd DC 0
VinCOA1 COA1 Gnd DC 0
VinCOA0 COA0 Gnd DC 0

VinCOB3 COB3 Gnd PULSE('SUPPLY' 0 0ns 100ps 100ps 40ns 80ns)
VinCOB2 COB2 Gnd PULSE('SUPPLY' 0 0ns 100ps 100ps 20ns 40ns)
VinCOB1 COB1 Gnd PULSE('SUPPLY' 0 0ns 100ps 100ps 10ns 20ns)
VinCOB0 COB0 Gnd PULSE('SUPPLY' 0 0ns 100ps 100ps 5ns 10ns)

M1000 COA1 COB1not EQ2 w_317_49# CMOSP w=20 l=2
+  ad=220 pd=62 as=440 ps=124
M1001 G G3 VDD VDD CMOSP w=20 l=2
+  ad=880 pd=248 as=7040 ps=1984
M1002 E1 a_416_140# Gnd Gnd CMOSN w=20 l=4
+  ad=220 pd=62 as=3740 ps=1054
M1003 G G2 VDD w_724_n227# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1004 a_352_n313# COA1 a_352_n353# Gnd CMOSN w=20 l=4
+  ad=440 pd=124 as=440 ps=124
M1005 COA0not COB0 EQ1 w_175_134# CMOSP w=20 l=2
+  ad=440 pd=124 as=440 ps=124
M1006 COB3not COB3 VDD VDD CMOSP w=20 l=2
+  ad=220 pd=62 as=0 ps=0
M1007 a_746_23# EQ3 a_746_n17# Gnd CMOSN w=20 l=4
+  ad=440 pd=124 as=440 ps=124
M1008 COA2not COA2 VDD VDD CMOSP w=20 l=2
+  ad=440 pd=124 as=0 ps=0
M1009 G3 COB0not VDD VDD CMOSP w=20 l=2
+  ad=1100 pd=310 as=0 ps=0
M1010 Gnd E1 L Gnd CMOSN w=20 l=4
+  ad=0 pd=0 as=440 ps=124
M1011 G1 COA2 VDD w_168_n228# CMOSP w=20 l=2
+  ad=660 pd=186 as=0 ps=0
M1012 COA1not COB1 EQ2 w_316_134# CMOSP w=20 l=2
+  ad=440 pd=124 as=0 ps=0
M1013 E1 a_416_140# VDD w_617_125# CMOSP w=20 l=2
+  ad=220 pd=62 as=0 ps=0
M1014 a_429_8# EQ4 Gnd Gnd CMOSN w=20 l=4
+  ad=440 pd=124 as=0 ps=0
M1015 a_352_n353# COB1not Gnd Gnd CMOSN w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1016 a_416_140# EQ3 VDD w_509_134# CMOSP w=20 l=2
+  ad=880 pd=248 as=0 ps=0
M1017 EQ3 COB2 COA2 Gnd CMOSN w=20 l=4
+  ad=420 pd=122 as=220 ps=62
M1018 G1 COB2not VDD VDD CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1019 G G0 VDD VDD CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1020 a_416_140# EQ1 VDD VDD CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1021 a_416_140# EQ1 a_429_88# Gnd CMOSN w=20 l=4
+  ad=220 pd=62 as=440 ps=124
M1022 COA2not COB2 EQ3 w_175_n47# CMOSP w=20 l=2
+  ad=0 pd=0 as=440 ps=124
M1023 EQ4 COB3not COA3not Gnd CMOSN w=20 l=4
+  ad=420 pd=122 as=440 ps=124
M1024 COA3 COB3not EQ4 w_317_n132# CMOSP w=20 l=2
+  ad=220 pd=62 as=440 ps=124
M1025 COB1not COB1 Gnd Gnd CMOSN w=20 l=4
+  ad=220 pd=62 as=0 ps=0
M1026 G3 COA0 VDD w_882_69# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1027 COA3not COB3 EQ4 w_316_n47# CMOSP w=20 l=2
+  ad=440 pd=124 as=0 ps=0
M1028 COA2 COB2not EQ3 w_176_n132# CMOSP w=20 l=2
+  ad=220 pd=62 as=0 ps=0
M1029 a_352_n273# EQ3 a_352_n313# Gnd CMOSN w=20 l=4
+  ad=440 pd=124 as=0 ps=0
M1030 a_429_48# EQ3 a_429_8# Gnd CMOSN w=20 l=4
+  ad=440 pd=124 as=0 ps=0
M1031 COB2not COB2 Gnd Gnd CMOSN w=20 l=4
+  ad=220 pd=62 as=0 ps=0
M1032 L G a_587_n123# w_581_n129# CMOSP w=20 l=2
+  ad=220 pd=62 as=440 ps=124
M1033 G1 EQ4 VDD VDD CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1034 COB0not COB0 VDD VDD CMOSP w=20 l=2
+  ad=220 pd=62 as=0 ps=0
M1035 a_416_140# EQ4 VDD VDD CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1036 a_644_n313# G2 a_644_n353# Gnd CMOSN w=20 l=4
+  ad=440 pd=124 as=440 ps=124
M1037 a_416_140# EQ2 VDD w_453_134# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1038 G3 EQ3 VDD w_770_69# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1039 a_429_88# EQ2 a_429_48# Gnd CMOSN w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1040 G3 EQ2 VDD w_826_69# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1041 COA3not COA3 VDD VDD CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1042 G2 EQ4 a_352_n273# Gnd CMOSN w=20 l=4
+  ad=220 pd=62 as=0 ps=0
M1043 COB2not COB2 VDD VDD CMOSP w=20 l=2
+  ad=220 pd=62 as=0 ps=0
M1044 a_644_n353# G3 Gnd Gnd CMOSN w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1045 a_459_n129# COB3not Gnd Gnd CMOSN w=20 l=4
+  ad=440 pd=124 as=0 ps=0
M1046 EQ2 COB1not COA1not Gnd CMOSN w=20 l=4
+  ad=420 pd=122 as=440 ps=124
M1047 COA3not COA3 Gnd Gnd CMOSN w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1048 G2 EQ3 VDD w_376_n227# CMOSP w=20 l=2
+  ad=880 pd=248 as=0 ps=0
M1049 a_144_n314# COB2not Gnd Gnd CMOSN w=20 l=4
+  ad=440 pd=124 as=0 ps=0
M1050 COA1not COA1 Gnd Gnd CMOSN w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1051 COB3not COB3 Gnd Gnd CMOSN w=20 l=4
+  ad=220 pd=62 as=0 ps=0
M1052 COA1not COA1 VDD VDD CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1053 G3 EQ4 VDD VDD CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1054 G0 COB3not VDD VDD CMOSP w=20 l=2
+  ad=440 pd=124 as=0 ps=0
M1055 a_644_n273# G1 a_644_n313# Gnd CMOSN w=20 l=4
+  ad=440 pd=124 as=0 ps=0
M1056 EQ1 COB0not COA0not Gnd CMOSN w=20 l=4
+  ad=420 pd=122 as=440 ps=124
M1057 G3 EQ4 a_746_23# Gnd CMOSN w=20 l=4
+  ad=220 pd=62 as=0 ps=0
M1058 G0 COA3 VDD VDD CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1059 EQ2 COB1 COA1 Gnd CMOSN w=20 l=4
+  ad=0 pd=0 as=220 ps=62
M1060 COA0not COA0 Gnd Gnd CMOSN w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1061 G0 COA3 a_459_n129# Gnd CMOSN w=20 l=4
+  ad=220 pd=62 as=0 ps=0
M1062 a_144_n274# COA2 a_144_n314# Gnd CMOSN w=20 l=4
+  ad=440 pd=124 as=0 ps=0
M1063 a_746_n96# COB0not Gnd Gnd CMOSN w=20 l=4
+  ad=440 pd=124 as=0 ps=0
M1064 EQ4 COB3 COA3 Gnd CMOSN w=20 l=4
+  ad=0 pd=0 as=220 ps=62
M1065 G2 EQ4 VDD VDD CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1066 COA0not COA0 VDD VDD CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1067 a_746_n17# EQ2 a_746_n57# Gnd CMOSN w=20 l=4
+  ad=0 pd=0 as=440 ps=124
M1068 G G0 a_644_n273# Gnd CMOSN w=20 l=4
+  ad=220 pd=62 as=0 ps=0
M1069 EQ1 COB0 COA0 Gnd CMOSN w=20 l=4
+  ad=0 pd=0 as=220 ps=62
M1070 COA0 COB0not EQ1 w_176_49# CMOSP w=20 l=2
+  ad=220 pd=62 as=0 ps=0
M1071 a_746_n57# COA0 a_746_n96# Gnd CMOSN w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1072 G2 COA1 VDD w_432_n227# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1073 COB1not COB1 VDD VDD CMOSP w=20 l=2
+  ad=220 pd=62 as=0 ps=0
M1074 COB0not COB0 Gnd Gnd CMOSN w=20 l=4
+  ad=220 pd=62 as=0 ps=0
M1075 EQ3 COB2not COA2not Gnd CMOSN w=20 l=4
+  ad=0 pd=0 as=440 ps=124
M1076 a_587_n123# E1 VDD VDD CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1077 COA2not COA2 Gnd Gnd CMOSN w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1078 Gnd G L Gnd CMOSN w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1079 G G1 VDD w_668_n227# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1080 G2 COB1not VDD VDD CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1081 G1 EQ4 a_144_n274# Gnd CMOSN w=20 l=4
+  ad=220 pd=62 as=0 ps=0
C0 w_509_134# a_416_140# 0.06fF
C1 COA3not Gnd 0.21fF
C2 G w_724_n227# 0.06fF
C3 EQ2 w_317_49# 0.09fF
C4 COB2 VDD 0.06fF
C5 EQ1 w_176_49# 0.09fF
C6 EQ2 w_316_134# 0.09fF
C7 a_352_n353# a_352_n313# 0.22fF
C8 a_746_n57# a_746_n96# 0.22fF
C9 E1 a_587_n123# 0.05fF
C10 w_176_49# COA0 0.06fF
C11 a_644_n353# Gnd 0.22fF
C12 COB0not VDD 0.40fF
C13 EQ4 w_317_n132# 0.09fF
C14 a_644_n273# G 0.21fF
C15 G2 EQ4 0.29fF
C16 COB1not w_317_49# 0.06fF
C17 G2 a_352_n273# 0.21fF
C18 COB3 w_316_n47# 0.06fF
C19 E1 w_617_125# 0.06fF
C20 COB1 COB1not 0.05fF
C21 VDD w_826_69# 0.09fF
C22 w_882_69# G3 0.06fF
C23 a_144_n314# a_144_n274# 0.21fF
C24 EQ3 w_176_n132# 0.09fF
C25 a_144_n314# Gnd 0.22fF
C26 G G3 0.16fF
C27 VDD w_724_n227# 0.09fF
C28 a_459_n129# Gnd 0.21fF
C29 COA3 G0 0.29fF
C30 EQ3 a_416_140# 0.16fF
C31 COA2not w_175_n47# 0.06fF
C32 w_509_134# VDD 0.09fF
C33 VDD COA1 0.06fF
C34 COA2not COB2not 0.01fF
C35 EQ1 a_416_140# 0.29fF
C36 L Gnd 0.41fF
C37 COB0not G3 0.16fF
C38 COA3not VDD 0.34fF
C39 COA1not w_316_134# 0.06fF
C40 G2 COB1not 0.16fF
C41 COA3 w_317_n132# 0.06fF
C42 w_882_69# COA0 0.06fF
C43 L w_581_n129# 0.06fF
C44 COB3not Gnd 0.21fF
C45 L G 0.25fF
C46 w_826_69# G3 0.06fF
C47 VDD G3 1.56fF
C48 a_746_n17# a_746_n57# 0.22fF
C49 COB3 COB3not 0.05fF
C50 EQ1 COB0not 0.25fF
C51 E1 Gnd 0.36fF
C52 G1 COB2not 0.16fF
C53 a_416_140# a_429_88# 0.21fF
C54 COA3 EQ4 0.68fF
C55 COB2not w_176_n132# 0.06fF
C56 COB2not Gnd 0.21fF
C57 COA3not w_316_n47# 0.06fF
C58 a_429_48# a_429_8# 0.22fF
C59 G G0 0.29fF
C60 VDD w_376_n227# 0.09fF
C61 EQ1 VDD 0.06fF
C62 EQ2 COB1not 0.25fF
C63 VDD COA0 0.06fF
C64 COA2 w_168_n228# 0.06fF
C65 EQ3 w_509_134# 0.06fF
C66 EQ1 w_175_134# 0.09fF
C67 COB2 w_175_n47# 0.06fF
C68 G2 G 0.16fF
C69 G1 EQ4 0.29fF
C70 COB2 COB2not 0.05fF
C71 COB3not VDD 0.40fF
C72 EQ2 w_453_134# 0.06fF
C73 COB1 VDD 0.06fF
C74 w_432_n227# VDD 0.09fF
C75 G1 COA2 0.16fF
C76 EQ4 a_416_140# 0.16fF
C77 COA2 w_176_n132# 0.06fF
C78 VDD G0 0.74fF
C79 EQ3 G3 0.16fF
C80 COA1not EQ2 0.68fF
C81 COA1 w_317_49# 0.06fF
C82 a_587_n123# w_581_n129# 0.09fF
C83 E1 VDD 0.27fF
C84 G1 w_668_n227# 0.06fF
C85 COA0not Gnd 0.21fF
C86 w_432_n227# COA1 0.06fF
C87 VDD COB2not 0.40fF
C88 COA0 G3 0.16fF
C89 COA3not COB3not 0.01fF
C90 EQ2 a_416_140# 0.16fF
C91 w_617_125# a_416_140# 0.06fF
C92 COA1not COB1not 0.01fF
C93 G2 VDD 1.22fF
C94 G2 w_724_n227# 0.06fF
C95 COA2not Gnd 0.21fF
C96 COB1not Gnd 0.21fF
C97 EQ3 w_376_n227# 0.06fF
C98 G w_668_n227# 0.06fF
C99 G1 w_168_n228# 0.06fF
C100 G2 COA1 0.16fF
C101 EQ1 COA0 0.68fF
C102 EQ4 VDD 0.26fF
C103 COA0not COB0not 0.01fF
C104 VDD a_587_n123# 0.34fF
C105 COA2 VDD 0.06fF
C106 w_453_134# a_416_140# 0.06fF
C107 VDD w_770_69# 0.09fF
C108 a_429_48# a_429_88# 0.21fF
C109 G1 a_144_n274# 0.21fF
C110 COA1not Gnd 0.21fF
C111 COB0not w_176_49# 0.06fF
C112 a_352_n273# a_352_n313# 0.21fF
C113 a_459_n129# G0 0.21fF
C114 EQ2 w_826_69# 0.06fF
C115 COA0not VDD 0.34fF
C116 w_617_125# VDD 0.06fF
C117 VDD w_668_n227# 0.09fF
C118 COA3not EQ4 0.68fF
C119 EQ3 w_175_n47# 0.09fF
C120 EQ3 COB2not 0.25fF
C121 COA0not w_175_134# 0.06fF
C122 G2 EQ3 0.16fF
C123 COB1 w_316_134# 0.06fF
C124 G1 G 0.16fF
C125 COA2not VDD 0.34fF
C126 VDD COB1not 0.40fF
C127 EQ4 w_316_n47# 0.09fF
C128 EQ2 COA1 0.68fF
C129 a_644_n273# a_644_n313# 0.21fF
C130 a_352_n353# Gnd 0.22fF
C131 EQ4 G3 0.29fF
C132 G Gnd 0.28fF
C133 G2 w_376_n227# 0.06fF
C134 COA3 VDD 0.13fF
C135 COB3not G0 0.16fF
C136 a_644_n313# a_644_n353# 0.22fF
C137 VDD w_168_n228# 0.09fF
C138 G w_581_n129# 0.06fF
C139 w_770_69# G3 0.06fF
C140 a_746_n96# Gnd 0.22fF
C141 COB0not COB0 0.05fF
C142 COB0not Gnd 0.21fF
C143 w_453_134# VDD 0.09fF
C144 EQ2 G3 0.16fF
C145 COB3not w_317_n132# 0.06fF
C146 COA1not VDD 0.34fF
C147 G2 w_432_n227# 0.06fF
C148 COA2 EQ3 0.68fF
C149 G1 VDD 0.95fF
C150 EQ3 w_770_69# 0.06fF
C151 COB0 VDD 0.06fF
C152 L a_587_n123# 0.27fF
C153 VDD Gnd 1.80fF
C154 a_429_8# Gnd 0.22fF
C155 a_746_23# G3 0.21fF
C156 VDD a_416_140# 1.22fF
C157 COB0 w_175_134# 0.06fF
C158 COB3 VDD 0.06fF
C159 a_746_23# a_746_n17# 0.21fF
C160 COA0not EQ1 0.68fF
C161 VDD w_882_69# 0.09fF
C162 COB3not EQ4 0.25fF
C163 G VDD 1.22fF
C164 COA2not EQ3 0.68fF
C165 Gnd Gnd 3.27fF
C166 G3 Gnd 1.66fF
C167 COB1not Gnd 0.99fF
C168 a_644_n353# Gnd 0.21fF
C169 a_352_n353# Gnd 0.21fF
C170 G2 Gnd 1.45fF
C171 COA1 Gnd 0.93fF
C172 COB2not Gnd 0.98fF
C173 a_644_n313# Gnd 0.22fF
C174 a_352_n313# Gnd 0.22fF
C175 a_144_n314# Gnd 0.22fF
C176 G1 Gnd 1.16fF
C177 EQ3 Gnd 1.65fF
C178 COA2 Gnd 0.86fF
C179 a_644_n273# Gnd 0.18fF
C180 a_352_n273# Gnd 0.18fF
C181 a_144_n274# Gnd 0.18fF
C182 G0 Gnd 0.70fF
C183 EQ4 Gnd 2.68fF
C184 G Gnd 1.42fF
C185 E1 Gnd 0.54fF
C186 COB3 Gnd 0.85fF
C187 COB3not Gnd 1.06fF
C188 COB2 Gnd 0.55fF
C189 COB0not Gnd 0.97fF
C190 L Gnd 0.17fF
C191 a_459_n129# Gnd 0.22fF
C192 COA3 Gnd 0.94fF
C193 COA3not Gnd 0.24fF
C194 COA2not Gnd 0.17fF
C195 a_746_n96# Gnd 0.21fF
C196 COA0 Gnd 0.72fF
C197 a_587_n123# Gnd 0.13fF
C198 a_746_n57# Gnd 0.21fF
C199 EQ2 Gnd 1.45fF
C200 a_746_n17# Gnd 0.22fF
C201 a_746_23# Gnd 0.18fF
C202 a_429_8# Gnd 0.21fF
C203 COB1 Gnd 0.81fF
C204 COB0 Gnd 0.63fF
C205 a_429_48# Gnd 0.22fF
C206 COA1not Gnd 0.22fF
C207 EQ1 Gnd 0.32fF
C208 COA0not Gnd 0.15fF
C209 a_429_88# Gnd 0.22fF
C210 a_416_140# Gnd 0.47fF
C211 w_724_n227# Gnd 1.16fF
C212 w_668_n227# Gnd 1.16fF
C213 VDD Gnd 21.24fF
C214 w_432_n227# Gnd 1.16fF
C215 w_376_n227# Gnd 1.16fF
C216 w_168_n228# Gnd 1.16fF
C217 w_581_n129# Gnd 1.16fF
C218 w_317_n132# Gnd 1.12fF
C219 w_176_n132# Gnd 1.16fF
C220 w_316_n47# Gnd 1.16fF
C221 w_175_n47# Gnd 0.67fF
C222 w_882_69# Gnd 1.16fF
C223 w_826_69# Gnd 1.16fF
C224 w_770_69# Gnd 1.16fF
C225 w_317_49# Gnd 1.16fF
C226 w_176_49# Gnd 0.61fF
C227 w_617_125# Gnd 1.16fF
C228 w_509_134# Gnd 1.16fF
C229 w_453_134# Gnd 1.16fF
C230 w_316_134# Gnd 1.16fF
C231 w_175_134# Gnd 0.67fF

.tran 1n 80ns
.control
run
set color0 = white
set color1 = black
plot v(L) v(E1)+2 v(G)+4
.endc
.end