Testing File for subcircuits

.include TSMC_180nm.txt

.include AND2.sub
.include AND3.sub
.include AND4.sub
.include NAND2.sub
.include NAND3.sub
.include NAND4.sub
.include NAND5.sub
.include NOR2.sub
.include NOT.sub
.include OR2.sub
.include XNOR2.sub
.include XOR2.sub

.include "FA.sub"

.include decoder.sub
.include Enable.sub
.include adder_subtractor.sub
.include comparator.sub
.include and_4bit.sub

.param SUPPLY = 1.8
.param LAMBDA = 0.18u

.param wn1 = {10*LAMBDA}
.param ln1 = {2*LAMBDA}
.param wn2 = {10*LAMBDA}
.param ln2 = {2*LAMBDA}
.param wn3 = {10*LAMBDA}
.param ln3 = {2*LAMBDA}
.param wn4 = {10*LAMBDA}
.param ln4 = {2*LAMBDA}
.param wn5 = {10*LAMBDA}
.param ln5 = {2*LAMBDA}

.param wp1 = wn1
.param lp1 = {LAMBDA}
.param wp2 = wn2
.param lp2 = {LAMBDA}
.param wp3 = wn3
.param lp3 = {LAMBDA}
.param wp4 = wn4
.param lp4 = {LAMBDA}
.param wp5 = wn5
.param lp5 = {LAMBDA}

.global GND

Vdd V GND 'SUPPLY'

* VA3 A3 GND PULSE(0 'SUPPLY' 0ns 100ps 100ps 80ns 160ns)
* VA2 A2 GND PULSE(0 'SUPPLY' 0ns 100ps 100ps 40ns 80ns)
* VA1 A1 GND PULSE(0 'SUPPLY' 0ns 100ps 100ps 20ns 40ns)
* VA0 A0 GND PULSE(0 'SUPPLY' 0ns 100ps 100ps 10ns 20ns)

VA3 A3 GND DC 0 ;'SUPPLY'
VA2 A2 GND DC 0 ;'SUPPLY'
VA1 A1 GND DC 0 ;'SUPPLY'
VA0 A0 GND DC 0 ;'SUPPLY'

VB3 B3 GND DC 'SUPPLY'
VB2 B2 GND DC 'SUPPLY'
VB1 B1 GND DC 'SUPPLY'
VB0 B0 GND DC 'SUPPLY'

VM M GND DC 0


Xtest A3 A2 A1 A0 B3 B2 B1 B0 M C S3 S2 S1 S0 V GND adder_subtractor

.tran 1n 160n

.control 
run
set color0 = rgb:f/f/e
set color1 = black
plot v(C)+8 v(S3)+6 v(S2)+4 v(S1)+2 v(S0)
.endc
.end