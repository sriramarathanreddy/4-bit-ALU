magic
tech scmos
timestamp 1701543619
<< nwell >>
rect 3355 -144 3391 -112
rect 3418 -144 3454 -112
rect 3496 -144 3532 -112
rect 3559 -144 3595 -112
rect 3640 -144 3676 -112
rect 3696 -144 3732 -112
rect 3752 -144 3788 -112
rect 3808 -144 3844 -112
rect 3860 -153 3896 -121
rect 3355 -226 3391 -194
rect 3419 -229 3455 -197
rect 3496 -226 3532 -194
rect 3560 -229 3596 -197
rect 3957 -209 3993 -177
rect 4013 -209 4049 -177
rect 4069 -209 4105 -177
rect 4125 -209 4161 -177
rect 4180 -209 4216 -177
rect 3355 -325 3391 -293
rect 3418 -325 3454 -293
rect 3496 -325 3532 -293
rect 3559 -325 3595 -293
rect 3670 -361 3706 -329
rect 3726 -361 3762 -329
rect 3824 -361 3860 -329
rect 3355 -407 3391 -375
rect 3419 -410 3455 -378
rect 3496 -407 3532 -375
rect 3560 -410 3596 -378
rect 3824 -407 3860 -375
rect 3355 -506 3391 -474
rect 3411 -506 3447 -474
rect 3467 -506 3503 -474
rect 3563 -505 3599 -473
rect 3619 -505 3655 -473
rect 3675 -505 3711 -473
rect 3731 -505 3767 -473
rect 3855 -505 3891 -473
rect 3911 -505 3947 -473
rect 3967 -505 4003 -473
rect 4023 -505 4059 -473
rect 4137 -583 4173 -551
rect 4193 -583 4229 -551
rect 4248 -592 4284 -560
<< ntransistor >>
rect 3371 -174 3375 -154
rect 3450 -183 3454 -163
rect 3512 -174 3516 -154
rect 3591 -183 3595 -163
rect 3683 -190 3687 -170
rect 3876 -183 3880 -163
rect 3683 -230 3687 -210
rect 3371 -256 3375 -236
rect 3451 -268 3455 -248
rect 3512 -256 3516 -236
rect 3592 -268 3596 -248
rect 3683 -270 3687 -250
rect 4000 -255 4004 -235
rect 3683 -309 3687 -289
rect 4000 -295 4004 -275
rect 4000 -335 4004 -315
rect 3371 -355 3375 -335
rect 3450 -364 3454 -344
rect 3512 -355 3516 -335
rect 3591 -364 3595 -344
rect 4000 -374 4004 -354
rect 3713 -407 3717 -387
rect 4000 -413 4004 -393
rect 3371 -437 3375 -417
rect 3451 -449 3455 -429
rect 3512 -437 3516 -417
rect 3592 -449 3596 -429
rect 3713 -447 3717 -427
rect 3830 -447 3834 -427
rect 3881 -447 3885 -427
rect 3398 -552 3402 -532
rect 3606 -551 3610 -531
rect 3898 -551 3902 -531
rect 3398 -592 3402 -572
rect 3606 -591 3610 -571
rect 3898 -591 3902 -571
rect 3398 -632 3402 -612
rect 3606 -631 3610 -611
rect 3898 -631 3902 -611
rect 4180 -629 4184 -609
rect 4264 -622 4268 -602
rect 3606 -670 3610 -650
rect 3898 -670 3902 -650
rect 4180 -669 4184 -649
<< ptransistor >>
rect 3372 -138 3374 -118
rect 3435 -138 3437 -118
rect 3513 -138 3515 -118
rect 3576 -138 3578 -118
rect 3657 -138 3659 -118
rect 3713 -138 3715 -118
rect 3769 -138 3771 -118
rect 3825 -138 3827 -118
rect 3877 -147 3879 -127
rect 3372 -220 3374 -200
rect 3436 -223 3438 -203
rect 3513 -220 3515 -200
rect 3974 -203 3976 -183
rect 4030 -203 4032 -183
rect 4086 -203 4088 -183
rect 4142 -203 4144 -183
rect 4197 -203 4199 -183
rect 3577 -223 3579 -203
rect 3372 -319 3374 -299
rect 3435 -319 3437 -299
rect 3513 -319 3515 -299
rect 3576 -319 3578 -299
rect 3687 -355 3689 -335
rect 3743 -355 3745 -335
rect 3841 -355 3843 -335
rect 3372 -401 3374 -381
rect 3436 -404 3438 -384
rect 3513 -401 3515 -381
rect 3577 -404 3579 -384
rect 3841 -401 3843 -381
rect 3372 -500 3374 -480
rect 3428 -500 3430 -480
rect 3484 -500 3486 -480
rect 3580 -499 3582 -479
rect 3636 -499 3638 -479
rect 3692 -499 3694 -479
rect 3748 -499 3750 -479
rect 3872 -499 3874 -479
rect 3928 -499 3930 -479
rect 3984 -499 3986 -479
rect 4040 -499 4042 -479
rect 4154 -577 4156 -557
rect 4210 -577 4212 -557
rect 4265 -586 4267 -566
<< ndiffusion >>
rect 3370 -174 3371 -154
rect 3375 -174 3376 -154
rect 3449 -183 3450 -163
rect 3454 -183 3455 -163
rect 3511 -174 3512 -154
rect 3516 -174 3517 -154
rect 3590 -183 3591 -163
rect 3595 -183 3596 -163
rect 3682 -190 3683 -170
rect 3687 -190 3688 -170
rect 3875 -183 3876 -163
rect 3880 -183 3881 -163
rect 3682 -230 3683 -210
rect 3687 -230 3688 -210
rect 3370 -256 3371 -236
rect 3375 -256 3376 -236
rect 3450 -268 3451 -248
rect 3455 -268 3456 -248
rect 3511 -256 3512 -236
rect 3516 -256 3517 -236
rect 3591 -268 3592 -248
rect 3596 -268 3597 -248
rect 3682 -270 3683 -250
rect 3687 -270 3688 -250
rect 3999 -255 4000 -235
rect 4004 -255 4005 -235
rect 3682 -309 3683 -289
rect 3687 -309 3688 -289
rect 3999 -295 4000 -275
rect 4004 -295 4005 -275
rect 3999 -335 4000 -315
rect 4004 -335 4005 -315
rect 3370 -355 3371 -335
rect 3375 -355 3376 -335
rect 3449 -364 3450 -344
rect 3454 -364 3455 -344
rect 3511 -355 3512 -335
rect 3516 -355 3517 -335
rect 3590 -364 3591 -344
rect 3595 -364 3596 -344
rect 3999 -374 4000 -354
rect 4004 -374 4005 -354
rect 3712 -407 3713 -387
rect 3717 -407 3718 -387
rect 3999 -413 4000 -393
rect 4004 -413 4005 -393
rect 3370 -437 3371 -417
rect 3375 -437 3376 -417
rect 3450 -449 3451 -429
rect 3455 -449 3456 -429
rect 3511 -437 3512 -417
rect 3516 -437 3517 -417
rect 3591 -449 3592 -429
rect 3596 -449 3597 -429
rect 3712 -447 3713 -427
rect 3717 -447 3718 -427
rect 3829 -447 3830 -427
rect 3834 -447 3835 -427
rect 3880 -447 3881 -427
rect 3885 -447 3886 -427
rect 3397 -552 3398 -532
rect 3402 -552 3403 -532
rect 3605 -551 3606 -531
rect 3610 -551 3611 -531
rect 3897 -551 3898 -531
rect 3902 -551 3903 -531
rect 3397 -592 3398 -572
rect 3402 -592 3403 -572
rect 3605 -591 3606 -571
rect 3610 -591 3611 -571
rect 3897 -591 3898 -571
rect 3902 -591 3903 -571
rect 3397 -632 3398 -612
rect 3402 -632 3403 -612
rect 3605 -631 3606 -611
rect 3610 -631 3611 -611
rect 3897 -631 3898 -611
rect 3902 -631 3903 -611
rect 4179 -629 4180 -609
rect 4184 -629 4185 -609
rect 4263 -622 4264 -602
rect 4268 -622 4269 -602
rect 3605 -670 3606 -650
rect 3610 -670 3611 -650
rect 3897 -670 3898 -650
rect 3902 -670 3903 -650
rect 4179 -669 4180 -649
rect 4184 -669 4185 -649
<< pdiffusion >>
rect 3371 -138 3372 -118
rect 3374 -138 3375 -118
rect 3434 -138 3435 -118
rect 3437 -138 3438 -118
rect 3512 -138 3513 -118
rect 3515 -138 3516 -118
rect 3575 -138 3576 -118
rect 3578 -138 3579 -118
rect 3656 -138 3657 -118
rect 3659 -138 3660 -118
rect 3712 -138 3713 -118
rect 3715 -138 3716 -118
rect 3768 -138 3769 -118
rect 3771 -138 3772 -118
rect 3824 -138 3825 -118
rect 3827 -138 3828 -118
rect 3876 -147 3877 -127
rect 3879 -147 3880 -127
rect 3371 -220 3372 -200
rect 3374 -220 3375 -200
rect 3435 -223 3436 -203
rect 3438 -223 3439 -203
rect 3512 -220 3513 -200
rect 3515 -220 3516 -200
rect 3973 -203 3974 -183
rect 3976 -203 3977 -183
rect 4029 -203 4030 -183
rect 4032 -203 4033 -183
rect 4085 -203 4086 -183
rect 4088 -203 4089 -183
rect 4141 -203 4142 -183
rect 4144 -203 4145 -183
rect 4196 -203 4197 -183
rect 4199 -203 4200 -183
rect 3576 -223 3577 -203
rect 3579 -223 3580 -203
rect 3371 -319 3372 -299
rect 3374 -319 3375 -299
rect 3434 -319 3435 -299
rect 3437 -319 3438 -299
rect 3512 -319 3513 -299
rect 3515 -319 3516 -299
rect 3575 -319 3576 -299
rect 3578 -319 3579 -299
rect 3686 -355 3687 -335
rect 3689 -355 3690 -335
rect 3742 -355 3743 -335
rect 3745 -355 3746 -335
rect 3840 -355 3841 -335
rect 3843 -355 3844 -335
rect 3371 -401 3372 -381
rect 3374 -401 3375 -381
rect 3435 -404 3436 -384
rect 3438 -404 3439 -384
rect 3512 -401 3513 -381
rect 3515 -401 3516 -381
rect 3576 -404 3577 -384
rect 3579 -404 3580 -384
rect 3840 -401 3841 -381
rect 3843 -401 3844 -381
rect 3371 -500 3372 -480
rect 3374 -500 3375 -480
rect 3427 -500 3428 -480
rect 3430 -500 3431 -480
rect 3483 -500 3484 -480
rect 3486 -500 3487 -480
rect 3579 -499 3580 -479
rect 3582 -499 3583 -479
rect 3635 -499 3636 -479
rect 3638 -499 3639 -479
rect 3691 -499 3692 -479
rect 3694 -499 3695 -479
rect 3747 -499 3748 -479
rect 3750 -499 3751 -479
rect 3871 -499 3872 -479
rect 3874 -499 3875 -479
rect 3927 -499 3928 -479
rect 3930 -499 3931 -479
rect 3983 -499 3984 -479
rect 3986 -499 3987 -479
rect 4039 -499 4040 -479
rect 4042 -499 4043 -479
rect 4153 -577 4154 -557
rect 4156 -577 4157 -557
rect 4209 -577 4210 -557
rect 4212 -577 4213 -557
rect 4264 -586 4265 -566
rect 4267 -586 4268 -566
<< ndcontact >>
rect 3360 -174 3370 -154
rect 3376 -174 3386 -154
rect 3439 -183 3449 -163
rect 3455 -183 3465 -163
rect 3501 -174 3511 -154
rect 3517 -174 3527 -154
rect 3580 -183 3590 -163
rect 3596 -183 3606 -163
rect 3672 -190 3682 -170
rect 3688 -190 3698 -170
rect 3865 -183 3875 -163
rect 3881 -183 3891 -163
rect 3672 -230 3682 -210
rect 3688 -230 3698 -210
rect 3360 -256 3370 -236
rect 3376 -256 3386 -236
rect 3440 -268 3450 -248
rect 3456 -268 3465 -248
rect 3501 -256 3511 -236
rect 3517 -256 3527 -236
rect 3581 -268 3591 -248
rect 3597 -268 3606 -248
rect 3672 -270 3682 -250
rect 3688 -270 3698 -250
rect 3989 -255 3999 -235
rect 4005 -255 4015 -235
rect 3672 -309 3682 -289
rect 3688 -309 3698 -289
rect 3989 -295 3999 -275
rect 4005 -295 4015 -275
rect 3989 -335 3999 -315
rect 4005 -335 4015 -315
rect 3360 -355 3370 -335
rect 3376 -355 3386 -335
rect 3439 -364 3449 -344
rect 3455 -364 3465 -344
rect 3501 -355 3511 -335
rect 3517 -355 3527 -335
rect 3580 -364 3590 -344
rect 3596 -364 3606 -344
rect 3989 -374 3999 -354
rect 4005 -374 4015 -354
rect 3702 -407 3712 -387
rect 3718 -407 3728 -387
rect 3989 -413 3999 -393
rect 4005 -413 4015 -393
rect 3360 -437 3370 -417
rect 3376 -437 3386 -417
rect 3440 -449 3450 -429
rect 3456 -449 3465 -429
rect 3501 -437 3511 -417
rect 3517 -437 3527 -417
rect 3581 -449 3591 -429
rect 3597 -449 3606 -429
rect 3702 -447 3712 -427
rect 3718 -447 3728 -427
rect 3819 -447 3829 -427
rect 3835 -447 3845 -427
rect 3870 -447 3880 -427
rect 3886 -447 3896 -427
rect 3387 -552 3397 -532
rect 3403 -552 3413 -532
rect 3595 -551 3605 -531
rect 3611 -551 3621 -531
rect 3887 -551 3897 -531
rect 3903 -551 3913 -531
rect 3387 -592 3397 -572
rect 3403 -592 3413 -572
rect 3595 -591 3605 -571
rect 3611 -591 3621 -571
rect 3887 -591 3897 -571
rect 3903 -591 3913 -571
rect 3387 -632 3397 -612
rect 3403 -632 3413 -612
rect 3595 -631 3605 -611
rect 3611 -631 3621 -611
rect 3887 -631 3897 -611
rect 3903 -631 3913 -611
rect 4169 -629 4179 -609
rect 4185 -629 4195 -609
rect 4253 -622 4263 -602
rect 4269 -622 4279 -602
rect 3595 -670 3605 -650
rect 3611 -670 3621 -650
rect 3887 -670 3897 -650
rect 3903 -670 3913 -650
rect 4169 -669 4179 -649
rect 4185 -669 4195 -649
<< pdcontact >>
rect 3361 -138 3371 -118
rect 3375 -138 3385 -118
rect 3424 -138 3434 -118
rect 3438 -138 3448 -118
rect 3502 -138 3512 -118
rect 3516 -138 3526 -118
rect 3565 -138 3575 -118
rect 3579 -138 3589 -118
rect 3646 -138 3656 -118
rect 3660 -138 3670 -118
rect 3702 -138 3712 -118
rect 3716 -138 3726 -118
rect 3758 -138 3768 -118
rect 3772 -138 3782 -118
rect 3814 -138 3824 -118
rect 3828 -138 3838 -118
rect 3866 -147 3876 -127
rect 3880 -147 3890 -127
rect 3361 -220 3371 -200
rect 3375 -220 3385 -200
rect 3425 -223 3435 -203
rect 3439 -223 3449 -203
rect 3502 -220 3512 -200
rect 3516 -220 3526 -200
rect 3963 -203 3973 -183
rect 3977 -203 3987 -183
rect 4019 -203 4029 -183
rect 4033 -203 4043 -183
rect 4075 -203 4085 -183
rect 4089 -203 4099 -183
rect 4131 -203 4141 -183
rect 4145 -203 4155 -183
rect 4186 -203 4196 -183
rect 4200 -203 4210 -183
rect 3566 -223 3576 -203
rect 3580 -223 3590 -203
rect 3361 -319 3371 -299
rect 3375 -319 3385 -299
rect 3424 -319 3434 -299
rect 3438 -319 3448 -299
rect 3502 -319 3512 -299
rect 3516 -319 3526 -299
rect 3565 -319 3575 -299
rect 3579 -319 3589 -299
rect 3676 -355 3686 -335
rect 3690 -355 3700 -335
rect 3732 -355 3742 -335
rect 3746 -355 3756 -335
rect 3830 -355 3840 -335
rect 3844 -355 3854 -335
rect 3361 -401 3371 -381
rect 3375 -401 3385 -381
rect 3425 -404 3435 -384
rect 3439 -404 3449 -384
rect 3502 -401 3512 -381
rect 3516 -401 3526 -381
rect 3566 -404 3576 -384
rect 3580 -404 3590 -384
rect 3830 -401 3840 -381
rect 3844 -401 3854 -381
rect 3361 -500 3371 -480
rect 3375 -500 3385 -480
rect 3417 -500 3427 -480
rect 3431 -500 3441 -480
rect 3473 -500 3483 -480
rect 3487 -500 3497 -480
rect 3569 -499 3579 -479
rect 3583 -499 3593 -479
rect 3625 -499 3635 -479
rect 3639 -499 3649 -479
rect 3681 -499 3691 -479
rect 3695 -499 3705 -479
rect 3737 -499 3747 -479
rect 3751 -499 3761 -479
rect 3861 -499 3871 -479
rect 3875 -499 3885 -479
rect 3917 -499 3927 -479
rect 3931 -499 3941 -479
rect 3973 -499 3983 -479
rect 3987 -499 3997 -479
rect 4029 -499 4039 -479
rect 4043 -499 4053 -479
rect 4143 -577 4153 -557
rect 4157 -577 4167 -557
rect 4199 -577 4209 -557
rect 4213 -577 4223 -557
rect 4254 -586 4264 -566
rect 4268 -586 4278 -566
<< psubstratepcontact >>
rect 3355 -184 3359 -180
rect 3387 -184 3391 -180
rect 3496 -184 3500 -180
rect 3528 -184 3532 -180
rect 3355 -266 3359 -262
rect 3387 -266 3391 -262
rect 3496 -266 3500 -262
rect 3528 -266 3532 -262
rect 3640 -318 3644 -314
rect 3840 -318 3844 -314
rect 3861 -318 3865 -314
rect 3893 -318 3897 -314
rect 3355 -365 3359 -361
rect 3387 -365 3391 -361
rect 3496 -365 3500 -361
rect 3528 -365 3532 -361
rect 3355 -447 3359 -443
rect 3387 -447 3391 -443
rect 3957 -422 3961 -418
rect 4212 -422 4216 -418
rect 3496 -447 3500 -443
rect 3528 -447 3532 -443
rect 3670 -457 3674 -453
rect 3758 -457 3762 -453
rect 3799 -461 3803 -457
rect 3892 -461 3896 -457
rect 3355 -641 3359 -637
rect 3499 -641 3503 -637
rect 3563 -679 3567 -675
rect 3763 -679 3767 -675
rect 3855 -679 3859 -675
rect 4055 -679 4059 -675
rect 4137 -679 4141 -675
rect 4225 -679 4229 -675
rect 4248 -679 4252 -675
rect 4280 -679 4284 -675
<< nsubstratencontact >>
rect 3355 -112 3359 -108
rect 3387 -112 3391 -108
rect 3496 -112 3500 -108
rect 3528 -112 3532 -108
rect 3640 -112 3644 -108
rect 3839 -112 3843 -108
rect 3861 -112 3865 -108
rect 3893 -112 3897 -108
rect 3957 -177 3961 -173
rect 4212 -177 4216 -173
rect 3355 -194 3359 -190
rect 3387 -194 3391 -190
rect 3496 -194 3500 -190
rect 3528 -194 3532 -190
rect 3355 -293 3359 -289
rect 3387 -293 3391 -289
rect 3496 -293 3500 -289
rect 3528 -293 3532 -289
rect 3670 -329 3674 -325
rect 3758 -329 3762 -325
rect 3824 -329 3828 -325
rect 3856 -329 3860 -325
rect 3355 -375 3359 -371
rect 3387 -375 3391 -371
rect 3496 -375 3500 -371
rect 3528 -375 3532 -371
rect 3355 -474 3359 -470
rect 3499 -474 3503 -470
rect 3563 -473 3567 -469
rect 3763 -473 3767 -469
rect 3855 -473 3859 -469
rect 4055 -473 4059 -469
rect 4137 -551 4141 -547
rect 4225 -551 4229 -547
rect 4248 -551 4252 -547
rect 4280 -551 4284 -547
<< polysilicon >>
rect 3372 -118 3374 -115
rect 3435 -118 3437 -115
rect 3513 -118 3515 -115
rect 3576 -118 3578 -115
rect 3657 -118 3659 -115
rect 3713 -118 3715 -115
rect 3769 -118 3771 -115
rect 3825 -118 3827 -115
rect 3877 -127 3879 -124
rect 3372 -147 3374 -138
rect 3435 -147 3437 -138
rect 3513 -147 3515 -138
rect 3576 -147 3578 -138
rect 3657 -147 3659 -138
rect 3713 -147 3715 -138
rect 3769 -147 3771 -138
rect 3825 -147 3827 -138
rect 3357 -149 3374 -147
rect 3357 -151 3375 -149
rect 3420 -151 3437 -147
rect 3498 -149 3515 -147
rect 3498 -151 3516 -149
rect 3561 -151 3578 -147
rect 3644 -151 3659 -147
rect 3700 -151 3715 -147
rect 3756 -151 3771 -147
rect 3812 -151 3827 -147
rect 3371 -154 3375 -151
rect 3512 -154 3516 -151
rect 3450 -163 3454 -160
rect 3371 -177 3375 -174
rect 3877 -156 3879 -147
rect 3862 -158 3879 -156
rect 3862 -160 3880 -158
rect 3591 -163 3595 -160
rect 3876 -163 3880 -160
rect 3512 -177 3516 -174
rect 3450 -186 3454 -183
rect 3672 -167 3687 -163
rect 3683 -170 3687 -167
rect 3591 -186 3595 -183
rect 3437 -190 3454 -186
rect 3578 -190 3595 -186
rect 3974 -183 3976 -180
rect 4030 -183 4032 -180
rect 4086 -183 4088 -180
rect 4142 -183 4144 -180
rect 4197 -183 4199 -180
rect 3876 -186 3880 -183
rect 3683 -193 3687 -190
rect 3372 -200 3374 -197
rect 3513 -200 3515 -197
rect 3436 -203 3438 -200
rect 3372 -229 3374 -220
rect 3577 -203 3579 -200
rect 3357 -231 3374 -229
rect 3357 -233 3375 -231
rect 3436 -232 3438 -223
rect 3513 -229 3515 -220
rect 3672 -207 3687 -203
rect 3683 -210 3687 -207
rect 3371 -236 3375 -233
rect 3421 -236 3438 -232
rect 3498 -231 3515 -229
rect 3498 -233 3516 -231
rect 3577 -232 3579 -223
rect 3974 -212 3976 -203
rect 4030 -212 4032 -203
rect 4086 -212 4088 -203
rect 4142 -212 4144 -203
rect 4197 -212 4199 -203
rect 3961 -216 3976 -212
rect 4017 -216 4032 -212
rect 4073 -216 4088 -212
rect 4129 -216 4144 -212
rect 4184 -216 4199 -212
rect 3512 -236 3516 -233
rect 3562 -236 3579 -232
rect 3683 -233 3687 -230
rect 3989 -232 4004 -228
rect 4000 -235 4004 -232
rect 3451 -248 3455 -245
rect 3371 -259 3375 -256
rect 3592 -248 3596 -245
rect 3672 -247 3687 -243
rect 3512 -259 3516 -256
rect 3683 -250 3687 -247
rect 3451 -271 3455 -268
rect 3592 -271 3596 -268
rect 4000 -258 4004 -255
rect 3438 -275 3455 -271
rect 3579 -275 3596 -271
rect 3683 -273 3687 -270
rect 3989 -272 4004 -268
rect 4000 -275 4004 -272
rect 3672 -286 3687 -282
rect 3683 -289 3687 -286
rect 3372 -299 3374 -296
rect 3435 -299 3437 -296
rect 3513 -299 3515 -296
rect 3576 -299 3578 -296
rect 4000 -298 4004 -295
rect 3683 -312 3687 -309
rect 3989 -312 4004 -308
rect 4000 -315 4004 -312
rect 3372 -328 3374 -319
rect 3435 -328 3437 -319
rect 3513 -328 3515 -319
rect 3576 -328 3578 -319
rect 3357 -330 3374 -328
rect 3357 -332 3375 -330
rect 3420 -332 3437 -328
rect 3498 -330 3515 -328
rect 3498 -332 3516 -330
rect 3561 -332 3578 -328
rect 3371 -335 3375 -332
rect 3512 -335 3516 -332
rect 3687 -335 3689 -332
rect 3743 -335 3745 -332
rect 3841 -335 3843 -332
rect 3450 -344 3454 -341
rect 3371 -358 3375 -355
rect 3591 -344 3595 -341
rect 3512 -358 3516 -355
rect 3450 -367 3454 -364
rect 4000 -338 4004 -335
rect 3989 -351 4004 -347
rect 4000 -354 4004 -351
rect 3687 -364 3689 -355
rect 3743 -364 3745 -355
rect 3841 -364 3843 -355
rect 3591 -367 3595 -364
rect 3437 -371 3454 -367
rect 3578 -371 3595 -367
rect 3674 -368 3689 -364
rect 3730 -368 3745 -364
rect 3828 -368 3843 -364
rect 4000 -377 4004 -374
rect 3372 -381 3374 -378
rect 3513 -381 3515 -378
rect 3436 -384 3438 -381
rect 3372 -410 3374 -401
rect 3577 -384 3579 -381
rect 3702 -384 3717 -380
rect 3841 -381 3843 -378
rect 3357 -412 3374 -410
rect 3357 -414 3375 -412
rect 3436 -413 3438 -404
rect 3513 -410 3515 -401
rect 3713 -387 3717 -384
rect 3371 -417 3375 -414
rect 3421 -417 3438 -413
rect 3498 -412 3515 -410
rect 3498 -414 3516 -412
rect 3577 -413 3579 -404
rect 3989 -390 4004 -386
rect 4000 -393 4004 -390
rect 3713 -410 3717 -407
rect 3841 -410 3843 -401
rect 3512 -417 3516 -414
rect 3562 -417 3579 -413
rect 3828 -414 3843 -410
rect 4000 -416 4004 -413
rect 3451 -429 3455 -426
rect 3371 -440 3375 -437
rect 3702 -424 3717 -420
rect 3592 -429 3596 -426
rect 3713 -427 3717 -424
rect 3830 -427 3834 -424
rect 3881 -427 3885 -424
rect 3512 -440 3516 -437
rect 3451 -452 3455 -449
rect 3592 -452 3596 -449
rect 3713 -450 3717 -447
rect 3830 -450 3834 -447
rect 3881 -450 3885 -447
rect 3438 -456 3455 -452
rect 3579 -456 3596 -452
rect 3817 -454 3834 -450
rect 3868 -454 3885 -450
rect 3372 -480 3374 -477
rect 3428 -480 3430 -477
rect 3484 -480 3486 -477
rect 3580 -479 3582 -476
rect 3636 -479 3638 -476
rect 3692 -479 3694 -476
rect 3748 -479 3750 -476
rect 3872 -479 3874 -476
rect 3928 -479 3930 -476
rect 3984 -479 3986 -476
rect 4040 -479 4042 -476
rect 3372 -509 3374 -500
rect 3428 -509 3430 -500
rect 3484 -509 3486 -500
rect 3580 -508 3582 -499
rect 3636 -508 3638 -499
rect 3692 -508 3694 -499
rect 3748 -508 3750 -499
rect 3872 -508 3874 -499
rect 3928 -508 3930 -499
rect 3984 -508 3986 -499
rect 4040 -508 4042 -499
rect 3359 -513 3374 -509
rect 3415 -513 3430 -509
rect 3471 -513 3486 -509
rect 3567 -512 3582 -508
rect 3623 -512 3638 -508
rect 3679 -512 3694 -508
rect 3735 -512 3750 -508
rect 3859 -512 3874 -508
rect 3915 -512 3930 -508
rect 3971 -512 3986 -508
rect 4027 -512 4042 -508
rect 3387 -529 3402 -525
rect 3595 -528 3610 -524
rect 3887 -528 3902 -524
rect 3398 -532 3402 -529
rect 3606 -531 3610 -528
rect 3898 -531 3902 -528
rect 3398 -555 3402 -552
rect 3606 -554 3610 -551
rect 3898 -554 3902 -551
rect 4154 -557 4156 -554
rect 4210 -557 4212 -554
rect 3387 -569 3402 -565
rect 3595 -568 3610 -564
rect 3887 -568 3902 -564
rect 3398 -572 3402 -569
rect 3606 -571 3610 -568
rect 3898 -571 3902 -568
rect 4265 -566 4267 -563
rect 4154 -586 4156 -577
rect 4210 -586 4212 -577
rect 4141 -590 4156 -586
rect 4197 -590 4212 -586
rect 3398 -595 3402 -592
rect 3606 -594 3610 -591
rect 3898 -594 3902 -591
rect 4265 -595 4267 -586
rect 4250 -597 4267 -595
rect 4250 -599 4268 -597
rect 4264 -602 4268 -599
rect 3387 -609 3402 -605
rect 3595 -608 3610 -604
rect 3887 -608 3902 -604
rect 4169 -606 4184 -602
rect 3398 -612 3402 -609
rect 3606 -611 3610 -608
rect 3898 -611 3902 -608
rect 4180 -609 4184 -606
rect 4264 -625 4268 -622
rect 3398 -635 3402 -632
rect 3606 -634 3610 -631
rect 3898 -634 3902 -631
rect 4180 -632 4184 -629
rect 3595 -647 3610 -643
rect 3887 -647 3902 -643
rect 4169 -646 4184 -642
rect 3606 -650 3610 -647
rect 3898 -650 3902 -647
rect 4180 -649 4184 -646
rect 3606 -673 3610 -670
rect 3898 -673 3902 -670
rect 4180 -672 4184 -669
<< polycontact >>
rect 3353 -151 3357 -147
rect 3416 -151 3420 -147
rect 3494 -151 3498 -147
rect 3557 -151 3561 -147
rect 3640 -151 3644 -147
rect 3696 -151 3700 -147
rect 3752 -151 3756 -147
rect 3808 -151 3812 -147
rect 3858 -160 3862 -156
rect 3668 -167 3672 -163
rect 3433 -190 3437 -186
rect 3574 -190 3578 -186
rect 3353 -233 3357 -229
rect 3668 -207 3672 -203
rect 3417 -236 3421 -232
rect 3494 -233 3498 -229
rect 3957 -216 3961 -212
rect 4013 -216 4017 -212
rect 4069 -216 4073 -212
rect 4125 -216 4129 -212
rect 4180 -216 4184 -212
rect 3558 -236 3562 -232
rect 3985 -232 3989 -228
rect 3668 -247 3672 -243
rect 3434 -275 3438 -271
rect 3575 -275 3579 -271
rect 3985 -272 3989 -268
rect 3668 -286 3672 -282
rect 3985 -312 3989 -308
rect 3353 -332 3357 -328
rect 3416 -332 3420 -328
rect 3494 -332 3498 -328
rect 3557 -332 3561 -328
rect 3985 -351 3989 -347
rect 3433 -371 3437 -367
rect 3574 -371 3578 -367
rect 3670 -368 3674 -364
rect 3726 -368 3730 -364
rect 3824 -368 3828 -364
rect 3698 -384 3702 -380
rect 3353 -414 3357 -410
rect 3417 -417 3421 -413
rect 3494 -414 3498 -410
rect 3985 -390 3989 -386
rect 3558 -417 3562 -413
rect 3824 -414 3828 -410
rect 3698 -424 3702 -420
rect 3434 -456 3438 -452
rect 3575 -456 3579 -452
rect 3813 -454 3817 -450
rect 3864 -454 3868 -450
rect 3355 -513 3359 -509
rect 3411 -513 3415 -509
rect 3467 -513 3471 -509
rect 3563 -512 3567 -508
rect 3619 -512 3623 -508
rect 3675 -512 3679 -508
rect 3731 -512 3735 -508
rect 3855 -512 3859 -508
rect 3911 -512 3915 -508
rect 3967 -512 3971 -508
rect 4023 -512 4027 -508
rect 3383 -529 3387 -525
rect 3591 -528 3595 -524
rect 3883 -528 3887 -524
rect 3383 -569 3387 -565
rect 3591 -568 3595 -564
rect 3883 -568 3887 -564
rect 4137 -590 4141 -586
rect 4193 -590 4197 -586
rect 4246 -599 4250 -595
rect 3383 -609 3387 -605
rect 3591 -608 3595 -604
rect 3883 -608 3887 -604
rect 4165 -606 4169 -602
rect 3591 -647 3595 -643
rect 3883 -647 3887 -643
rect 4165 -646 4169 -642
<< metal1 >>
rect 3359 -112 3387 -108
rect 3418 -112 3465 -108
rect 3500 -112 3528 -108
rect 3559 -112 3606 -108
rect 3644 -112 3839 -108
rect 3843 -112 3861 -108
rect 3865 -112 3893 -108
rect 3361 -118 3371 -112
rect 3424 -118 3434 -112
rect 3376 -147 3385 -138
rect 3339 -151 3353 -147
rect 3376 -151 3399 -147
rect 3402 -151 3416 -147
rect 3376 -154 3385 -151
rect 3439 -163 3448 -138
rect 3455 -163 3465 -112
rect 3502 -118 3512 -112
rect 3565 -118 3575 -112
rect 3517 -147 3526 -138
rect 3480 -151 3494 -147
rect 3517 -151 3540 -147
rect 3543 -151 3557 -147
rect 3517 -154 3526 -151
rect 3360 -180 3370 -174
rect 3359 -184 3387 -180
rect 3580 -163 3589 -138
rect 3596 -163 3606 -112
rect 3646 -118 3656 -112
rect 3702 -118 3712 -112
rect 3758 -118 3768 -112
rect 3814 -118 3824 -112
rect 3625 -151 3640 -147
rect 3660 -156 3670 -138
rect 3681 -151 3696 -147
rect 3716 -156 3726 -138
rect 3737 -151 3752 -147
rect 3772 -156 3782 -138
rect 3793 -151 3808 -147
rect 3828 -156 3838 -138
rect 3866 -127 3876 -112
rect 3881 -156 3890 -147
rect 3640 -160 3858 -156
rect 3881 -160 3904 -156
rect 3501 -180 3511 -174
rect 3500 -184 3528 -180
rect 3653 -167 3668 -163
rect 3688 -170 3698 -160
rect 3881 -163 3890 -160
rect 3419 -190 3433 -186
rect 3560 -190 3574 -186
rect 3961 -177 4212 -173
rect 3963 -183 3973 -177
rect 4019 -183 4029 -177
rect 4075 -183 4085 -177
rect 4131 -183 4141 -177
rect 4186 -183 4196 -177
rect 3359 -194 3387 -190
rect 3361 -200 3371 -194
rect 3419 -197 3465 -193
rect 3500 -194 3528 -190
rect 3376 -229 3385 -220
rect 3425 -203 3435 -197
rect 3339 -233 3353 -229
rect 3376 -233 3399 -229
rect 3376 -236 3385 -233
rect 3403 -236 3417 -232
rect 3440 -248 3449 -223
rect 3456 -248 3465 -197
rect 3502 -200 3512 -194
rect 3560 -197 3606 -193
rect 3517 -229 3526 -220
rect 3566 -203 3576 -197
rect 3480 -233 3494 -229
rect 3517 -233 3540 -229
rect 3517 -236 3526 -233
rect 3544 -236 3558 -232
rect 3360 -262 3370 -256
rect 3359 -266 3387 -262
rect 3581 -248 3590 -223
rect 3597 -248 3606 -197
rect 3672 -196 3682 -190
rect 3672 -200 3698 -196
rect 3653 -207 3668 -203
rect 3688 -210 3698 -200
rect 3672 -236 3682 -230
rect 3672 -240 3698 -236
rect 3653 -247 3668 -243
rect 3501 -262 3511 -256
rect 3500 -266 3528 -262
rect 3688 -250 3698 -240
rect 3420 -275 3434 -271
rect 3561 -275 3575 -271
rect 3672 -275 3682 -270
rect 3672 -279 3698 -275
rect 3653 -286 3668 -282
rect 3688 -289 3698 -279
rect 3359 -293 3387 -289
rect 3418 -293 3465 -289
rect 3500 -293 3528 -289
rect 3559 -293 3606 -289
rect 3361 -299 3371 -293
rect 3424 -299 3434 -293
rect 3376 -328 3385 -319
rect 3339 -332 3353 -328
rect 3376 -332 3399 -328
rect 3402 -332 3416 -328
rect 3376 -335 3385 -332
rect 3439 -344 3448 -319
rect 3455 -344 3465 -293
rect 3502 -299 3512 -293
rect 3565 -299 3575 -293
rect 3517 -328 3526 -319
rect 3480 -332 3494 -328
rect 3517 -332 3540 -328
rect 3543 -332 3557 -328
rect 3517 -335 3526 -332
rect 3360 -361 3370 -355
rect 3359 -365 3387 -361
rect 3580 -344 3589 -319
rect 3596 -344 3606 -293
rect 3672 -314 3682 -309
rect 3865 -314 3875 -183
rect 3942 -216 3957 -212
rect 3977 -221 3987 -203
rect 3998 -216 4013 -212
rect 4033 -221 4043 -203
rect 4054 -216 4069 -212
rect 4089 -221 4099 -203
rect 4110 -216 4125 -212
rect 4145 -221 4155 -203
rect 4165 -216 4180 -212
rect 4200 -221 4210 -203
rect 3957 -225 4216 -221
rect 3970 -232 3985 -228
rect 4005 -235 4015 -225
rect 3989 -261 3999 -255
rect 3989 -265 4015 -261
rect 3970 -272 3985 -268
rect 4005 -275 4015 -265
rect 3989 -301 3999 -295
rect 3989 -305 4015 -301
rect 3970 -312 3985 -308
rect 3644 -318 3840 -314
rect 3844 -318 3861 -314
rect 3865 -318 3893 -314
rect 4005 -315 4015 -305
rect 3674 -329 3758 -325
rect 3799 -329 3824 -325
rect 3828 -329 3856 -325
rect 3860 -329 3896 -325
rect 3501 -361 3511 -355
rect 3500 -365 3528 -361
rect 3676 -335 3686 -329
rect 3732 -335 3742 -329
rect 3830 -335 3840 -329
rect 3989 -340 3999 -335
rect 3989 -344 4015 -340
rect 3970 -351 3985 -347
rect 4005 -354 4015 -344
rect 3419 -371 3433 -367
rect 3560 -371 3574 -367
rect 3655 -368 3670 -364
rect 3359 -375 3387 -371
rect 3361 -381 3371 -375
rect 3419 -378 3465 -374
rect 3500 -375 3528 -371
rect 3690 -373 3700 -355
rect 3711 -368 3726 -364
rect 3746 -373 3756 -355
rect 3810 -368 3824 -364
rect 3844 -371 3854 -355
rect 3376 -410 3385 -401
rect 3425 -384 3435 -378
rect 3339 -414 3353 -410
rect 3376 -414 3399 -410
rect 3376 -417 3385 -414
rect 3403 -417 3417 -413
rect 3440 -429 3449 -404
rect 3456 -429 3465 -378
rect 3502 -381 3512 -375
rect 3560 -378 3606 -374
rect 3670 -377 3762 -373
rect 3824 -375 3860 -371
rect 3517 -410 3526 -401
rect 3566 -384 3576 -378
rect 3480 -414 3494 -410
rect 3517 -414 3540 -410
rect 3517 -417 3526 -414
rect 3544 -417 3558 -413
rect 3360 -443 3370 -437
rect 3359 -447 3387 -443
rect 3581 -429 3590 -404
rect 3597 -429 3606 -378
rect 3683 -384 3698 -380
rect 3718 -387 3728 -377
rect 3830 -381 3840 -375
rect 3989 -379 3999 -374
rect 3989 -383 4015 -379
rect 3970 -390 3985 -386
rect 4005 -393 4015 -383
rect 3702 -413 3712 -407
rect 3702 -417 3728 -413
rect 3810 -414 3824 -410
rect 3844 -417 3854 -401
rect 3683 -424 3698 -420
rect 3718 -427 3728 -417
rect 3799 -421 3896 -417
rect 3989 -418 3999 -413
rect 3501 -443 3511 -437
rect 3500 -447 3528 -443
rect 3819 -427 3829 -421
rect 3870 -427 3880 -421
rect 3961 -422 4212 -418
rect 3420 -456 3434 -452
rect 3561 -456 3575 -452
rect 3702 -453 3712 -447
rect 3674 -457 3758 -453
rect 3799 -454 3813 -450
rect 3835 -457 3845 -447
rect 3850 -454 3864 -450
rect 3886 -457 3896 -447
rect 3803 -461 3892 -457
rect 3359 -474 3499 -470
rect 3567 -473 3763 -469
rect 3859 -473 4055 -469
rect 3361 -480 3371 -474
rect 3417 -480 3427 -474
rect 3473 -480 3483 -474
rect 3569 -479 3579 -473
rect 3625 -479 3635 -473
rect 3681 -479 3691 -473
rect 3737 -479 3747 -473
rect 3861 -479 3871 -473
rect 3917 -479 3927 -473
rect 3973 -479 3983 -473
rect 4029 -479 4039 -473
rect 3340 -513 3355 -509
rect 3375 -518 3385 -500
rect 3396 -513 3411 -509
rect 3431 -518 3441 -500
rect 3452 -513 3467 -509
rect 3487 -518 3497 -500
rect 3548 -512 3563 -508
rect 3583 -517 3593 -499
rect 3604 -512 3619 -508
rect 3639 -517 3649 -499
rect 3660 -512 3675 -508
rect 3695 -517 3705 -499
rect 3716 -512 3731 -508
rect 3751 -517 3761 -499
rect 3840 -512 3855 -508
rect 3875 -517 3885 -499
rect 3896 -512 3911 -508
rect 3931 -517 3941 -499
rect 3952 -512 3967 -508
rect 3987 -517 3997 -499
rect 4008 -512 4023 -508
rect 4043 -517 4053 -499
rect 3355 -522 3503 -518
rect 3563 -521 3767 -517
rect 3855 -521 4059 -517
rect 3368 -529 3383 -525
rect 3403 -532 3413 -522
rect 3576 -528 3591 -524
rect 3611 -531 3621 -521
rect 3868 -528 3883 -524
rect 3903 -531 3913 -521
rect 4141 -551 4225 -547
rect 4229 -551 4248 -547
rect 4252 -551 4280 -547
rect 3387 -558 3397 -552
rect 3595 -557 3605 -551
rect 3887 -557 3897 -551
rect 4143 -557 4153 -551
rect 4199 -557 4209 -551
rect 3387 -562 3413 -558
rect 3595 -561 3621 -557
rect 3887 -561 3913 -557
rect 3368 -569 3383 -565
rect 3403 -572 3413 -562
rect 3576 -568 3591 -564
rect 3611 -571 3621 -561
rect 3868 -568 3883 -564
rect 3903 -571 3913 -561
rect 4122 -590 4137 -586
rect 3387 -598 3397 -592
rect 3595 -597 3605 -591
rect 3887 -597 3897 -591
rect 4157 -595 4167 -577
rect 4178 -590 4193 -586
rect 4213 -595 4223 -577
rect 4254 -566 4264 -551
rect 4269 -595 4278 -586
rect 3387 -602 3413 -598
rect 3595 -601 3621 -597
rect 3887 -601 3913 -597
rect 4137 -599 4246 -595
rect 4269 -599 4292 -595
rect 3368 -609 3383 -605
rect 3403 -612 3413 -602
rect 3576 -608 3591 -604
rect 3611 -611 3621 -601
rect 3868 -608 3883 -604
rect 3903 -611 3913 -601
rect 4150 -606 4165 -602
rect 4185 -609 4195 -599
rect 4269 -602 4278 -599
rect 3387 -637 3397 -632
rect 3595 -636 3605 -631
rect 3887 -636 3897 -631
rect 4169 -635 4179 -629
rect 3359 -641 3499 -637
rect 3595 -640 3621 -636
rect 3887 -640 3913 -636
rect 4169 -639 4195 -635
rect 3576 -647 3591 -643
rect 3611 -650 3621 -640
rect 3868 -647 3883 -643
rect 3903 -650 3913 -640
rect 4150 -646 4165 -642
rect 4185 -649 4195 -639
rect 3595 -675 3605 -670
rect 3887 -675 3897 -670
rect 4169 -675 4179 -669
rect 4253 -675 4263 -622
rect 3567 -679 3763 -675
rect 3859 -679 4055 -675
rect 4141 -679 4225 -675
rect 4229 -679 4248 -675
rect 4252 -679 4280 -675
<< labels >>
rlabel metal1 3355 -474 3503 -470 5 VDD
rlabel metal1 3355 -641 3503 -637 1 Gnd
rlabel metal1 3563 -679 3767 -675 1 Gnd
rlabel metal1 3563 -473 3767 -469 5 VDD
rlabel metal1 3855 -679 4059 -675 1 Gnd
rlabel metal1 3855 -473 4059 -469 5 VDD
rlabel metal1 3355 -112 3391 -108 5 VDD
rlabel metal1 3355 -184 3391 -180 1 Gnd
rlabel metal1 3355 -194 3391 -190 5 VDD
rlabel metal1 3355 -266 3391 -262 1 Gnd
rlabel metal1 3496 -112 3532 -108 5 VDD
rlabel metal1 3496 -184 3532 -180 1 Gnd
rlabel metal1 3496 -194 3532 -190 5 VDD
rlabel metal1 3496 -266 3532 -262 1 Gnd
rlabel metal1 3355 -293 3391 -289 5 VDD
rlabel metal1 3355 -365 3391 -361 1 Gnd
rlabel metal1 3355 -375 3391 -371 5 VDD
rlabel metal1 3355 -447 3391 -443 1 Gnd
rlabel metal1 3496 -293 3532 -289 5 VDD
rlabel metal1 3496 -365 3532 -361 1 Gnd
rlabel metal1 3496 -375 3532 -371 5 VDD
rlabel metal1 3496 -447 3532 -443 1 Gnd
rlabel metal1 3339 -151 3357 -147 1 COB0
rlabel metal1 3381 -151 3399 -147 1 COB0not
rlabel metal1 3339 -233 3357 -229 1 COA0
rlabel metal1 3381 -233 3399 -229 1 COA0not
rlabel metal1 3480 -151 3498 -147 1 COB1
rlabel metal1 3522 -151 3540 -147 1 COB1not
rlabel metal1 3480 -233 3498 -229 1 COA1
rlabel metal1 3522 -233 3540 -229 1 COA1not
rlabel metal1 3339 -332 3357 -328 1 COB2
rlabel metal1 3381 -332 3399 -328 1 COB2not
rlabel metal1 3339 -414 3357 -410 1 COA2
rlabel metal1 3381 -414 3399 -410 1 COA2not
rlabel metal1 3480 -332 3498 -328 1 COB3
rlabel metal1 3522 -332 3540 -328 1 COB3not
rlabel metal1 3480 -414 3498 -410 1 COA3
rlabel metal1 3522 -414 3540 -410 1 COA3not
rlabel metal1 3402 -151 3420 -147 1 COB0
rlabel metal1 3419 -190 3437 -186 1 COB0not
rlabel metal1 3403 -236 3421 -232 1 COB0not
rlabel metal1 3420 -275 3438 -271 1 COB0
rlabel metal1 3439 -163 3448 -138 1 COA0not
rlabel metal1 3440 -248 3449 -223 1 COA0
rlabel metal1 3455 -163 3465 -108 1 EQ1
rlabel metal1 3456 -248 3465 -193 1 EQ1
rlabel metal1 3543 -151 3561 -147 1 COB1
rlabel metal1 3561 -275 3579 -271 1 COB1
rlabel metal1 3560 -190 3578 -186 1 COB1not
rlabel metal1 3544 -236 3562 -232 1 COB1not
rlabel metal1 3580 -163 3589 -138 1 COA1not
rlabel metal1 3581 -248 3590 -223 1 COA1
rlabel metal1 3597 -248 3606 -193 1 EQ2
rlabel metal1 3596 -163 3606 -108 1 EQ2
rlabel metal1 3402 -332 3420 -328 1 COB2
rlabel metal1 3420 -456 3438 -452 1 COB2
rlabel metal1 3419 -371 3437 -367 1 COB2not
rlabel metal1 3403 -417 3421 -413 1 COB2not
rlabel metal1 3440 -429 3449 -404 1 COA2
rlabel metal1 3439 -344 3448 -319 1 COA2not
rlabel metal1 3456 -429 3465 -374 1 EQ3
rlabel metal1 3455 -344 3465 -289 1 EQ3
rlabel metal1 3596 -344 3606 -289 1 EQ4
rlabel metal1 3597 -429 3606 -374 1 EQ4
rlabel metal1 3580 -344 3589 -319 1 COA3not
rlabel metal1 3581 -429 3590 -404 1 COA3
rlabel metal1 3543 -332 3561 -328 1 COB3
rlabel metal1 3561 -456 3579 -452 1 COB3
rlabel metal1 3560 -371 3578 -367 1 COB3not
rlabel metal1 3544 -417 3562 -413 1 COB3not
rlabel metal1 3640 -112 3897 -108 5 VDD
rlabel metal1 3640 -318 3897 -314 1 Gnd
rlabel metal1 3625 -151 3644 -147 1 EQ1
rlabel metal1 3653 -167 3672 -163 1 EQ1
rlabel metal1 3681 -151 3700 -147 1 EQ2
rlabel metal1 3653 -207 3672 -203 1 EQ2
rlabel metal1 3737 -151 3756 -147 1 EQ3
rlabel metal1 3653 -247 3672 -243 1 EQ3
rlabel metal1 3653 -286 3672 -282 1 EQ4
rlabel metal1 3793 -151 3812 -147 1 EQ4
rlabel metal1 3885 -160 3904 -156 1 E1
rlabel metal1 3670 -457 3762 -453 1 Gnd
rlabel metal1 3670 -329 3762 -325 5 VDD
rlabel metal1 3799 -329 3896 -325 5 VDD
rlabel metal1 3799 -461 3896 -457 1 Gnd
rlabel metal1 3655 -368 3674 -364 1 COA3
rlabel metal1 3683 -384 3702 -380 1 COA3
rlabel metal1 3711 -368 3730 -364 1 COB3not
rlabel metal1 3683 -424 3702 -420 1 COB3not
rlabel metal1 3670 -377 3762 -373 1 G0
rlabel metal1 3810 -368 3828 -364 1 E1
rlabel metal1 3799 -454 3817 -450 1 E1
rlabel metal1 3810 -414 3828 -410 1 G
rlabel metal1 3850 -454 3868 -450 1 G
rlabel metal1 3799 -421 3896 -417 1 L
rlabel metal1 3957 -422 4216 -418 1 Gnd
rlabel metal1 3957 -177 4216 -173 5 VDD
rlabel metal1 3396 -513 3415 -509 1 COA2
rlabel metal1 3368 -569 3387 -565 1 COA2
rlabel metal1 3452 -513 3471 -509 1 COB2not
rlabel metal1 3368 -609 3387 -605 1 COB2not
rlabel metal1 3355 -522 3503 -518 1 G1
rlabel metal1 3563 -521 3767 -517 1 G2
rlabel metal1 3548 -512 3567 -508 1 EQ4
rlabel metal1 3340 -513 3359 -509 1 EQ4
rlabel metal1 3368 -529 3387 -525 1 EQ4
rlabel metal1 3576 -528 3595 -524 1 EQ4
rlabel metal1 3604 -512 3623 -508 1 EQ3
rlabel metal1 3576 -568 3595 -564 1 EQ3
rlabel metal1 3660 -512 3679 -508 1 COA1
rlabel metal1 3576 -608 3595 -604 1 COA1
rlabel metal1 3716 -512 3735 -508 1 COB1not
rlabel metal1 3576 -647 3595 -643 1 COB1not
rlabel metal1 3942 -216 3961 -212 1 EQ4
rlabel metal1 3970 -232 3989 -228 1 EQ4
rlabel metal1 3998 -216 4017 -212 1 EQ3
rlabel metal1 3970 -272 3989 -268 1 EQ3
rlabel metal1 4054 -216 4073 -212 1 EQ2
rlabel metal1 3970 -312 3989 -308 1 EQ2
rlabel metal1 4110 -216 4129 -212 1 COA0
rlabel metal1 3970 -351 3989 -347 1 COA0
rlabel metal1 4165 -216 4184 -212 1 COB0not
rlabel metal1 3970 -390 3989 -386 1 COB0not
rlabel metal1 3957 -225 4216 -221 1 G3
rlabel metal1 3840 -512 3859 -508 1 G0
rlabel metal1 3868 -528 3887 -524 1 G0
rlabel metal1 3896 -512 3915 -508 1 G1
rlabel metal1 3868 -568 3887 -564 1 G1
rlabel metal1 3952 -512 3971 -508 1 G2
rlabel metal1 3868 -608 3887 -604 1 G2
rlabel metal1 4008 -512 4027 -508 1 G3
rlabel metal1 3868 -647 3887 -643 1 G3
rlabel metal1 3855 -521 4059 -517 1 G
rlabel metal1 4137 -679 4284 -675 1 Gnd
rlabel metal1 4137 -551 4284 -547 5 VDD
rlabel metal1 4122 -590 4141 -586 1 E1
rlabel metal1 4150 -606 4169 -602 1 E1
rlabel metal1 4178 -590 4197 -586 1 D2
rlabel metal1 4150 -646 4169 -642 1 D2
rlabel metal1 4273 -599 4292 -595 1 E
<< end >>
