* SPICE3 file created from and_4bit.ext - technology: scmos

.include TSMC_180nm.txt
.param SUPPLY = 1.8
.global Gnd
Vdd VDD Gnd 'SUPPLY'
.option scale=0.09u

VinANA3 ANA3 Gnd DC 'SUPPLY'
VinANA2 ANA2 Gnd DC 0
VinANA1 ANA1 Gnd DC 'SUPPLY'
VinANA0 ANA0 Gnd DC 'SUPPLY'

VinANB3 ANB3 Gnd DC 'SUPPLY'
VinANB2 ANB2 Gnd DC 'SUPPLY'
VinANB1 ANB1 Gnd DC 0
VinANB0 ANB0 Gnd DC 'SUPPLY'

M1000 OUT_AND0 a_411_103# VDD w_503_88# CMOSP w=20 l=2
+  ad=220 pd=62 as=2640 ps=744
M1001 OUT_AND1 a_609_103# VDD w_701_88# CMOSP w=20 l=2
+  ad=220 pd=62 as=0 ps=0
M1002 OUT_AND2 a_807_103# VDD w_899_88# CMOSP w=20 l=2
+  ad=220 pd=62 as=0 ps=0
M1003 OUT_AND0 a_411_103# Gnd Gnd CMOSN w=20 l=4
+  ad=220 pd=62 as=1760 ps=496
M1004 OUT_AND1 a_609_103# Gnd Gnd CMOSN w=20 l=4
+  ad=220 pd=62 as=0 ps=0
M1005 OUT_AND3 a_1005_103# VDD w_1097_88# CMOSP w=20 l=2
+  ad=220 pd=62 as=0 ps=0
M1006 OUT_AND2 a_807_103# Gnd Gnd CMOSN w=20 l=4
+  ad=220 pd=62 as=0 ps=0
M1007 a_411_103# ANA0 a_424_51# Gnd CMOSN w=20 l=4
+  ad=220 pd=62 as=440 ps=124
M1008 OUT_AND3 a_1005_103# Gnd Gnd CMOSN w=20 l=4
+  ad=220 pd=62 as=0 ps=0
M1009 a_609_103# ANA1 a_622_51# Gnd CMOSN w=20 l=4
+  ad=220 pd=62 as=440 ps=124
M1010 a_807_103# ANA2 a_820_51# Gnd CMOSN w=20 l=4
+  ad=220 pd=62 as=440 ps=124
M1011 a_411_103# ANA0 VDD VDD CMOSP w=20 l=2
+  ad=440 pd=124 as=0 ps=0
M1012 a_609_103# ANA1 VDD VDD CMOSP w=20 l=2
+  ad=440 pd=124 as=0 ps=0
M1013 a_1005_103# ANB3 VDD VDD CMOSP w=20 l=2
+  ad=440 pd=124 as=0 ps=0
M1014 a_807_103# ANA2 VDD VDD CMOSP w=20 l=2
+  ad=440 pd=124 as=0 ps=0
M1015 a_1005_103# ANA3 VDD VDD CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1016 a_424_51# ANB0 Gnd Gnd CMOSN w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1017 a_1005_103# ANA3 a_1018_51# Gnd CMOSN w=20 l=4
+  ad=220 pd=62 as=440 ps=124
M1018 a_622_51# ANB1 Gnd Gnd CMOSN w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1019 a_820_51# ANB2 Gnd Gnd CMOSN w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1020 a_411_103# ANB0 VDD VDD CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1021 a_609_103# ANB1 VDD VDD CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1022 a_807_103# ANB2 VDD VDD CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1023 a_1018_51# ANB3 Gnd Gnd CMOSN w=20 l=4
+  ad=0 pd=0 as=0 ps=0
C0 ANB0 a_411_103# 0.10fF
C1 Gnd a_820_51# 0.21fF
C2 OUT_AND2 w_899_88# 0.06fF
C3 a_807_103# a_820_51# 0.21fF
C4 VDD w_899_88# 0.06fF
C5 w_1097_88# a_1005_103# 0.06fF
C6 a_424_51# Gnd 0.21fF
C7 OUT_AND2 VDD 0.21fF
C8 a_411_103# ANA0 0.47fF
C9 OUT_AND1 w_701_88# 0.06fF
C10 OUT_AND1 Gnd 0.14fF
C11 a_609_103# a_622_51# 0.21fF
C12 VDD OUT_AND3 0.21fF
C13 a_609_103# VDD 0.67fF
C14 OUT_AND0 w_503_88# 0.06fF
C15 ANB3 VDD 0.06fF
C16 ANB2 a_807_103# 0.10fF
C17 ANA2 VDD 0.06fF
C18 ANB0 VDD 0.06fF
C19 VDD ANA0 0.06fF
C20 Gnd a_622_51# 0.21fF
C21 a_807_103# w_899_88# 0.06fF
C22 VDD w_701_88# 0.06fF
C23 OUT_AND2 Gnd 0.14fF
C24 OUT_AND3 Gnd 0.14fF
C25 a_807_103# VDD 0.67fF
C26 a_609_103# w_701_88# 0.06fF
C27 ANB3 a_1018_51# 0.19fF
C28 VDD a_1005_103# 0.67fF
C29 OUT_AND0 VDD 0.21fF
C30 a_411_103# w_503_88# 0.06fF
C31 a_411_103# a_424_51# 0.21fF
C32 ANB2 a_820_51# 0.19fF
C33 ANA3 VDD 0.06fF
C34 ANB1 a_622_51# 0.19fF
C35 ANB3 a_1005_103# 0.10fF
C36 ANA2 a_807_103# 0.47fF
C37 ANB1 VDD 0.06fF
C38 ANB1 a_609_103# 0.10fF
C39 Gnd a_1018_51# 0.21fF
C40 VDD w_1097_88# 0.06fF
C41 w_1097_88# OUT_AND3 0.06fF
C42 a_1005_103# a_1018_51# 0.21fF
C43 VDD w_503_88# 0.06fF
C44 OUT_AND1 VDD 0.21fF
C45 OUT_AND0 Gnd 0.14fF
C46 a_411_103# VDD 0.67fF
C47 ANB2 VDD 0.06fF
C48 ANA3 a_1005_103# 0.47fF
C49 ANA1 VDD 0.06fF
C50 ANB0 a_424_51# 0.19fF
C51 ANA1 a_609_103# 0.47fF
C52 a_1018_51# Gnd 0.20fF
C53 a_820_51# Gnd 0.20fF
C54 a_622_51# Gnd 0.20fF
C55 Gnd Gnd 0.32fF
C56 a_424_51# Gnd 0.20fF
C57 OUT_AND3 Gnd 0.13fF
C58 a_1005_103# Gnd 0.78fF
C59 OUT_AND2 Gnd 0.13fF
C60 a_807_103# Gnd 0.78fF
C61 OUT_AND1 Gnd 0.13fF
C62 a_609_103# Gnd 0.78fF
C63 OUT_AND0 Gnd 0.13fF
C64 a_411_103# Gnd 0.78fF
C65 ANB3 Gnd 0.99fF
C66 ANA3 Gnd 0.54fF
C67 ANB2 Gnd 0.99fF
C68 ANA2 Gnd 0.57fF
C69 ANB1 Gnd 0.99fF
C70 ANA1 Gnd 0.59fF
C71 ANB0 Gnd 0.99fF
C72 ANA0 Gnd 0.62fF
C73 w_1097_88# Gnd 1.16fF
C74 w_899_88# Gnd 0.22fF
C75 w_701_88# Gnd 0.22fF
C76 w_503_88# Gnd 0.22fF
C77 VDD Gnd 11.46fF

.tran 1n 10n
.control
run
set color0 = white
set color1 = black
plot v(OUT_AND0) v(OUT_AND1)+2 v(OUT_AND2)+4 v(OUT_AND3)+6
.endc
.end