magic
tech scmos
timestamp 1701499843
<< nwell >>
rect 201 136 237 168
rect 257 136 293 168
rect 313 136 349 168
rect 365 127 401 159
<< ntransistor >>
rect 244 90 248 110
rect 244 50 248 70
rect 381 97 385 117
rect 244 10 248 30
<< ptransistor >>
rect 218 142 220 162
rect 274 142 276 162
rect 330 142 332 162
rect 382 133 384 153
<< ndiffusion >>
rect 243 90 244 110
rect 248 90 249 110
rect 243 50 244 70
rect 248 50 249 70
rect 380 97 381 117
rect 385 97 386 117
rect 243 10 244 30
rect 248 10 249 30
<< pdiffusion >>
rect 217 142 218 162
rect 220 142 221 162
rect 273 142 274 162
rect 276 142 277 162
rect 329 142 330 162
rect 332 142 333 162
rect 381 133 382 153
rect 384 133 385 153
<< ndcontact >>
rect 233 90 243 110
rect 249 90 259 110
rect 233 50 243 70
rect 249 50 259 70
rect 370 97 380 117
rect 386 97 396 117
rect 233 10 243 30
rect 249 10 259 30
<< pdcontact >>
rect 207 142 217 162
rect 221 142 231 162
rect 263 142 273 162
rect 277 142 287 162
rect 319 142 329 162
rect 333 142 343 162
rect 371 133 381 153
rect 385 133 395 153
<< psubstratepcontact >>
rect 201 1 205 5
rect 345 1 349 5
rect 365 1 369 5
rect 397 1 401 5
<< nsubstratencontact >>
rect 201 168 205 172
rect 345 168 349 172
rect 365 168 369 172
rect 397 168 401 172
<< polysilicon >>
rect 218 162 220 165
rect 274 162 276 165
rect 330 162 332 165
rect 382 153 384 156
rect 218 133 220 142
rect 274 133 276 142
rect 330 133 332 142
rect 205 129 220 133
rect 261 129 276 133
rect 317 129 332 133
rect 233 113 248 117
rect 244 110 248 113
rect 244 87 248 90
rect 272 77 276 129
rect 233 73 276 77
rect 244 70 248 73
rect 244 47 248 50
rect 328 37 332 129
rect 382 124 384 133
rect 367 122 384 124
rect 367 120 385 122
rect 381 117 385 120
rect 381 94 385 97
rect 233 33 332 37
rect 244 30 248 33
rect 244 7 248 10
<< polycontact >>
rect 201 129 205 133
rect 229 113 233 117
rect 229 73 233 77
rect 363 120 367 124
rect 229 33 233 37
<< metal1 >>
rect 205 168 345 172
rect 349 168 365 172
rect 369 168 397 172
rect 207 162 217 168
rect 263 162 273 168
rect 319 162 329 168
rect 186 129 201 133
rect 186 117 190 129
rect 221 124 231 142
rect 277 124 287 142
rect 333 124 343 142
rect 371 153 381 168
rect 386 124 395 133
rect 201 120 363 124
rect 386 120 409 124
rect 186 113 229 117
rect 249 110 259 120
rect 386 117 395 120
rect 233 84 243 90
rect 233 80 259 84
rect 214 73 229 77
rect 249 70 259 80
rect 233 44 243 50
rect 233 40 259 44
rect 214 33 229 37
rect 249 30 259 40
rect 233 5 243 10
rect 370 5 380 97
rect 205 1 345 5
rect 349 1 365 5
rect 369 1 397 5
<< labels >>
rlabel metal1 186 129 205 133 1 A
rlabel metal1 214 73 233 77 1 B
rlabel metal1 214 33 233 37 1 C
rlabel metal1 201 168 401 172 5 VDD
rlabel metal1 201 1 401 5 1 Gnd
rlabel metal1 390 120 409 124 1 OUT
<< end >>
