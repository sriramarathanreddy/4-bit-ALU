magic
tech scmos
timestamp 1701541558
<< nwell >>
rect 1667 8393 1902 8425
rect 1667 8388 1903 8393
rect 1668 8376 1903 8388
rect 1936 8305 1989 8330
rect 1936 8304 1982 8305
rect 4666 7932 4900 7964
rect 3710 7903 3820 7917
rect 3904 7910 3939 7911
rect 2668 7867 2771 7881
rect 2986 7872 3089 7886
rect 1777 7836 1887 7850
rect 1971 7843 2006 7844
rect 1778 7806 1887 7836
rect 1894 7809 2006 7843
rect 2176 7835 2286 7849
rect 2668 7846 2772 7867
rect 2986 7851 3090 7872
rect 3304 7870 3407 7884
rect 3711 7873 3820 7903
rect 3827 7876 3939 7910
rect 4180 7909 4290 7923
rect 4374 7916 4409 7917
rect 3904 7875 3939 7876
rect 3788 7872 3820 7873
rect 3962 7872 4015 7898
rect 4181 7879 4290 7909
rect 4297 7882 4409 7916
rect 4666 7916 4901 7932
rect 4666 7915 4841 7916
rect 4852 7915 4901 7916
rect 4374 7881 4409 7882
rect 4258 7878 4290 7879
rect 4432 7878 4485 7904
rect 2370 7842 2405 7843
rect 1971 7808 2006 7809
rect 1820 7805 1843 7806
rect 1855 7805 1887 7806
rect 2029 7805 2082 7831
rect 2177 7805 2286 7835
rect 2293 7808 2405 7842
rect 2370 7807 2405 7808
rect 2219 7804 2242 7805
rect 2254 7804 2286 7805
rect 2428 7804 2481 7830
rect 2668 7826 2769 7846
rect 2986 7831 3087 7851
rect 3304 7849 3408 7870
rect 3304 7829 3405 7849
rect 4934 7843 4988 7869
rect 2662 7697 2697 7718
rect 2980 7702 3015 7723
rect 3298 7700 3333 7721
rect 3068 7661 3106 7662
rect 2750 7656 2788 7657
rect 2616 7582 2670 7608
rect 2683 7605 2788 7656
rect 2934 7587 2988 7613
rect 3001 7610 3106 7661
rect 3386 7659 3424 7660
rect 3252 7585 3306 7611
rect 3319 7608 3424 7659
rect 2971 7127 3074 7141
rect 2617 7112 2720 7126
rect 1776 7081 1886 7095
rect 1970 7088 2005 7089
rect 1777 7051 1886 7081
rect 1893 7054 2005 7088
rect 2177 7086 2287 7100
rect 2371 7093 2406 7094
rect 1970 7053 2005 7054
rect 1819 7050 1842 7051
rect 1854 7050 1886 7051
rect 2028 7050 2081 7076
rect 2178 7056 2287 7086
rect 2294 7059 2406 7093
rect 2617 7091 2721 7112
rect 2971 7106 3075 7127
rect 3314 7125 3417 7139
rect 3713 7131 3823 7145
rect 3907 7138 3942 7139
rect 2371 7058 2406 7059
rect 2220 7055 2243 7056
rect 2255 7055 2287 7056
rect 2429 7055 2482 7081
rect 2617 7071 2718 7091
rect 2971 7086 3072 7106
rect 3314 7104 3418 7125
rect 3314 7084 3415 7104
rect 3714 7101 3823 7131
rect 3830 7104 3942 7138
rect 4183 7137 4293 7151
rect 4377 7144 4412 7145
rect 3907 7103 3942 7104
rect 3791 7100 3823 7101
rect 3965 7100 4018 7126
rect 4184 7107 4293 7137
rect 4300 7110 4412 7144
rect 4377 7109 4412 7110
rect 4261 7106 4293 7107
rect 4435 7106 4488 7132
rect 4666 7130 4900 7162
rect 4666 7114 4901 7130
rect 4666 7113 4841 7114
rect 4852 7113 4901 7114
rect 4934 7041 4988 7067
rect 2611 6942 2646 6963
rect 2965 6957 3000 6978
rect 3308 6955 3343 6976
rect 3053 6916 3091 6917
rect 2699 6901 2737 6902
rect 2565 6827 2619 6853
rect 2632 6850 2737 6901
rect 2919 6842 2973 6868
rect 2986 6865 3091 6916
rect 3396 6914 3434 6915
rect 3262 6840 3316 6866
rect 3329 6863 3434 6914
rect 2641 6221 2744 6235
rect 2947 6221 3050 6235
rect 3312 6234 3415 6248
rect 1777 6190 1887 6204
rect 1971 6197 2006 6198
rect 1778 6160 1887 6190
rect 1894 6163 2006 6197
rect 2178 6195 2288 6209
rect 2372 6202 2407 6203
rect 1971 6162 2006 6163
rect 1820 6159 1843 6160
rect 1855 6159 1887 6160
rect 2029 6159 2082 6185
rect 2179 6165 2288 6195
rect 2295 6168 2407 6202
rect 2641 6200 2745 6221
rect 2947 6200 3051 6221
rect 3312 6213 3416 6234
rect 2372 6167 2407 6168
rect 2221 6164 2244 6165
rect 2256 6164 2288 6165
rect 2430 6164 2483 6190
rect 2641 6180 2742 6200
rect 2947 6180 3048 6200
rect 3312 6193 3413 6213
rect 3713 6183 3823 6197
rect 3907 6190 3942 6191
rect 3714 6153 3823 6183
rect 3830 6156 3942 6190
rect 4183 6189 4293 6203
rect 4377 6196 4412 6197
rect 3907 6155 3942 6156
rect 3791 6152 3823 6153
rect 3965 6152 4018 6178
rect 4184 6159 4293 6189
rect 4300 6162 4412 6196
rect 4377 6161 4412 6162
rect 4261 6158 4293 6159
rect 4435 6158 4488 6184
rect 4666 6179 4900 6211
rect 4666 6163 4901 6179
rect 4666 6162 4841 6163
rect 4852 6162 4901 6163
rect 4934 6090 4988 6116
rect 2635 6051 2670 6072
rect 2941 6051 2976 6072
rect 3306 6064 3341 6085
rect 3394 6023 3432 6024
rect 2723 6010 2761 6011
rect 3029 6010 3067 6011
rect 2589 5936 2643 5962
rect 2656 5959 2761 6010
rect 2895 5936 2949 5962
rect 2962 5959 3067 6010
rect 3260 5949 3314 5975
rect 3327 5972 3432 6023
rect 3713 5520 3823 5534
rect 3907 5527 3942 5528
rect 3714 5490 3823 5520
rect 3830 5493 3942 5527
rect 4183 5526 4293 5540
rect 4377 5533 4412 5534
rect 3907 5492 3942 5493
rect 3791 5489 3823 5490
rect 3965 5489 4018 5515
rect 4184 5496 4293 5526
rect 4300 5499 4412 5533
rect 4377 5498 4412 5499
rect 4261 5495 4293 5496
rect 4435 5495 4488 5521
rect 4666 5515 4900 5547
rect 4666 5499 4901 5515
rect 4666 5498 4841 5499
rect 4852 5498 4901 5499
rect 2617 5441 2720 5455
rect 2959 5451 3062 5465
rect 3350 5460 3453 5474
rect 1775 5410 1885 5424
rect 1969 5417 2004 5418
rect 1776 5380 1885 5410
rect 1892 5383 2004 5417
rect 2176 5415 2286 5429
rect 2370 5422 2405 5423
rect 1969 5382 2004 5383
rect 1818 5379 1841 5380
rect 1853 5379 1885 5380
rect 2027 5379 2080 5405
rect 2177 5385 2286 5415
rect 2293 5388 2405 5422
rect 2617 5420 2721 5441
rect 2959 5430 3063 5451
rect 3350 5439 3454 5460
rect 2370 5387 2405 5388
rect 2219 5384 2242 5385
rect 2254 5384 2286 5385
rect 2428 5384 2481 5410
rect 2617 5400 2718 5420
rect 2959 5410 3060 5430
rect 3350 5419 3451 5439
rect 4934 5426 4988 5452
rect 2611 5271 2646 5292
rect 2953 5281 2988 5302
rect 3344 5290 3379 5311
rect 3432 5249 3470 5250
rect 3041 5240 3079 5241
rect 2699 5230 2737 5231
rect 2565 5156 2619 5182
rect 2632 5179 2737 5230
rect 2907 5166 2961 5192
rect 2974 5189 3079 5240
rect 3298 5175 3352 5201
rect 3365 5198 3470 5249
<< ntransistor >>
rect 1965 8280 1970 8285
rect 1708 8250 1719 8259
rect 1799 8250 1810 8259
rect 2057 7781 2060 7786
rect 1829 7678 1836 7689
rect 1938 7679 1945 7689
rect 2456 7780 2459 7785
rect 2708 7769 2715 7779
rect 3026 7774 3033 7784
rect 3344 7772 3351 7782
rect 3990 7848 3995 7853
rect 4460 7854 4465 7859
rect 4963 7819 4968 7824
rect 4706 7789 4717 7798
rect 4797 7789 4808 7798
rect 3756 7746 3769 7762
rect 3872 7749 3885 7765
rect 4226 7752 4239 7768
rect 4342 7755 4355 7771
rect 2228 7677 2235 7688
rect 2338 7677 2346 7688
rect 2991 7688 2993 7692
rect 2673 7683 2675 7687
rect 3309 7686 3311 7690
rect 2645 7558 2650 7563
rect 2963 7563 2968 7568
rect 2727 7548 2734 7558
rect 3045 7553 3052 7563
rect 3281 7561 3286 7566
rect 3363 7551 3370 7561
rect 2056 7026 2059 7031
rect 2457 7031 2460 7036
rect 3011 7029 3018 7039
rect 3354 7027 3361 7037
rect 2657 7014 2664 7024
rect 3993 7076 3998 7081
rect 4463 7082 4468 7087
rect 3759 6974 3772 6990
rect 3875 6977 3888 6993
rect 4229 6980 4242 6996
rect 4345 6983 4358 6999
rect 4963 7017 4968 7022
rect 4706 6987 4717 6996
rect 4797 6987 4808 6996
rect 1828 6923 1835 6934
rect 1938 6923 1945 6934
rect 2229 6928 2236 6939
rect 2339 6928 2347 6939
rect 2976 6943 2978 6947
rect 3319 6941 3321 6945
rect 2622 6928 2624 6932
rect 2948 6818 2953 6823
rect 2594 6803 2599 6808
rect 3030 6808 3037 6818
rect 3291 6816 3296 6821
rect 2676 6793 2683 6803
rect 3373 6806 3380 6816
rect 2057 6135 2060 6140
rect 1829 6032 1836 6043
rect 1938 6031 1945 6043
rect 2458 6140 2461 6145
rect 3352 6136 3359 6146
rect 2681 6123 2688 6133
rect 2987 6123 2994 6133
rect 2230 6037 2237 6048
rect 2338 6036 2346 6048
rect 3317 6050 3319 6054
rect 3993 6128 3998 6133
rect 4463 6134 4468 6139
rect 2646 6037 2648 6041
rect 2952 6037 2954 6041
rect 3759 6026 3772 6042
rect 3875 6029 3888 6045
rect 4229 6032 4242 6048
rect 4345 6035 4358 6051
rect 4963 6066 4968 6071
rect 4706 6036 4717 6045
rect 4797 6036 4808 6045
rect 2618 5912 2623 5917
rect 3289 5925 3294 5930
rect 2924 5912 2929 5917
rect 3371 5915 3378 5925
rect 2700 5902 2707 5912
rect 3006 5902 3013 5912
rect 2055 5355 2058 5360
rect 3993 5465 3998 5470
rect 4463 5471 4468 5476
rect 2456 5360 2459 5365
rect 2999 5353 3006 5363
rect 3390 5362 3397 5372
rect 3759 5363 3772 5379
rect 3875 5366 3888 5382
rect 4229 5369 4243 5385
rect 4345 5372 4358 5388
rect 4963 5402 4968 5407
rect 4706 5372 4717 5381
rect 4797 5372 4808 5381
rect 2657 5343 2664 5353
rect 1827 5252 1834 5263
rect 1937 5252 1946 5263
rect 2228 5257 2235 5268
rect 2338 5258 2344 5268
rect 3355 5276 3357 5280
rect 2964 5267 2966 5271
rect 2622 5257 2624 5261
rect 3327 5151 3332 5156
rect 2936 5142 2941 5147
rect 2594 5132 2599 5137
rect 3018 5132 3025 5142
rect 3409 5141 3416 5151
rect 2676 5122 2683 5132
<< ptransistor >>
rect 1708 8395 1719 8404
rect 1799 8395 1810 8404
rect 1965 8314 1970 8319
rect 1829 7815 1836 7831
rect 1939 7818 1946 7834
rect 2057 7815 2060 7820
rect 2228 7814 2235 7830
rect 2338 7817 2345 7833
rect 2705 7833 2713 7843
rect 3023 7838 3031 7848
rect 3756 7882 3769 7898
rect 3872 7885 3889 7901
rect 4226 7888 4239 7904
rect 4706 7934 4717 7943
rect 4797 7934 4808 7943
rect 4341 7891 4357 7907
rect 3341 7836 3349 7846
rect 2456 7814 2459 7819
rect 3990 7882 3995 7887
rect 4460 7888 4465 7893
rect 4963 7853 4968 7858
rect 2991 7708 2993 7712
rect 2673 7703 2675 7707
rect 3309 7706 3311 7710
rect 1828 7060 1835 7076
rect 1938 7063 1945 7079
rect 2229 7065 2236 7081
rect 2723 7612 2736 7622
rect 3041 7617 3054 7627
rect 3359 7615 3372 7625
rect 2963 7597 2968 7602
rect 2645 7592 2650 7597
rect 3281 7595 3286 7600
rect 2339 7068 2346 7084
rect 3008 7093 3016 7103
rect 3758 7110 3772 7126
rect 3875 7113 3888 7129
rect 4229 7116 4242 7132
rect 4345 7119 4358 7135
rect 4706 7132 4717 7141
rect 4797 7132 4808 7141
rect 3351 7091 3359 7101
rect 2654 7078 2662 7088
rect 2056 7060 2059 7065
rect 2457 7065 2460 7070
rect 3993 7110 3998 7115
rect 4463 7116 4468 7121
rect 4963 7051 4968 7056
rect 2976 6963 2978 6967
rect 2622 6948 2624 6952
rect 3319 6961 3321 6965
rect 1829 6169 1836 6185
rect 1938 6172 1945 6188
rect 2230 6174 2237 6190
rect 3026 6872 3039 6882
rect 3369 6870 3382 6880
rect 2672 6857 2685 6867
rect 2948 6852 2953 6857
rect 2594 6837 2599 6842
rect 3291 6850 3296 6855
rect 2340 6177 2347 6193
rect 3349 6200 3357 6210
rect 2678 6187 2686 6197
rect 2984 6187 2992 6197
rect 2057 6169 2060 6174
rect 2458 6174 2461 6179
rect 3759 6162 3772 6178
rect 3875 6165 3891 6181
rect 4229 6168 4242 6184
rect 4344 6171 4360 6187
rect 4706 6181 4717 6190
rect 4797 6181 4808 6190
rect 3317 6070 3319 6074
rect 2646 6057 2648 6061
rect 2952 6057 2954 6061
rect 1827 5389 1834 5405
rect 3993 6162 3998 6167
rect 4463 6168 4468 6173
rect 1937 5392 1945 5408
rect 2228 5394 2235 5410
rect 4963 6100 4968 6105
rect 3367 5979 3380 5989
rect 2696 5966 2709 5976
rect 3002 5966 3015 5976
rect 3289 5959 3294 5964
rect 2618 5946 2623 5951
rect 2924 5946 2929 5951
rect 3759 5499 3772 5515
rect 3873 5502 3888 5518
rect 4229 5505 4242 5521
rect 4345 5508 4361 5524
rect 4706 5517 4717 5526
rect 4797 5517 4808 5526
rect 2338 5397 2345 5413
rect 2996 5417 3004 5427
rect 3387 5426 3395 5436
rect 2654 5407 2662 5417
rect 2055 5389 2058 5394
rect 2456 5394 2459 5399
rect 3993 5499 3998 5504
rect 4463 5505 4468 5510
rect 4963 5436 4968 5441
rect 3355 5296 3357 5300
rect 2964 5287 2966 5291
rect 2622 5277 2624 5281
rect 3014 5196 3027 5206
rect 3405 5205 3418 5215
rect 2672 5186 2685 5196
rect 3327 5185 3332 5190
rect 2936 5176 2941 5181
rect 2594 5166 2599 5171
<< ndiffusion >>
rect 1960 8280 1965 8285
rect 1970 8280 1977 8285
rect 1676 8257 1708 8259
rect 1676 8250 1680 8257
rect 1691 8250 1708 8257
rect 1719 8258 1749 8259
rect 1719 8251 1734 8258
rect 1745 8251 1749 8258
rect 1719 8250 1749 8251
rect 1753 8257 1799 8259
rect 1753 8250 1757 8257
rect 1768 8250 1799 8257
rect 1810 8257 1850 8259
rect 1810 8250 1826 8257
rect 1837 8250 1850 8257
rect 2051 7781 2057 7786
rect 2060 7781 2069 7786
rect 1769 7688 1829 7689
rect 1796 7678 1829 7688
rect 1836 7679 1938 7689
rect 1945 7682 1988 7689
rect 1993 7682 1994 7689
rect 2451 7780 2456 7785
rect 2459 7780 2468 7785
rect 2677 7771 2681 7779
rect 2688 7771 2708 7779
rect 2677 7769 2708 7771
rect 2715 7771 2746 7779
rect 2753 7771 2757 7779
rect 2995 7776 2999 7784
rect 3006 7776 3026 7784
rect 2995 7774 3026 7776
rect 3033 7776 3064 7784
rect 3071 7776 3075 7784
rect 3033 7774 3075 7776
rect 3313 7774 3317 7782
rect 3324 7774 3344 7782
rect 2715 7769 2757 7771
rect 3313 7772 3344 7774
rect 3351 7774 3382 7782
rect 3389 7774 3393 7782
rect 3351 7772 3393 7774
rect 3985 7848 3990 7853
rect 3995 7848 4002 7853
rect 4455 7854 4460 7859
rect 4465 7854 4472 7859
rect 4958 7819 4963 7824
rect 4968 7819 4975 7824
rect 4674 7796 4706 7798
rect 4674 7789 4678 7796
rect 4689 7789 4706 7796
rect 4717 7797 4747 7798
rect 4717 7790 4732 7797
rect 4743 7790 4747 7797
rect 4717 7789 4747 7790
rect 4751 7796 4797 7798
rect 4751 7789 4755 7796
rect 4766 7789 4797 7796
rect 4808 7796 4848 7798
rect 4808 7789 4824 7796
rect 4835 7789 4848 7796
rect 4337 7770 4342 7771
rect 4289 7768 4342 7770
rect 3867 7764 3872 7765
rect 3819 7762 3872 7764
rect 3721 7757 3756 7762
rect 3721 7747 3729 7757
rect 3740 7747 3756 7757
rect 3721 7746 3756 7747
rect 3769 7749 3872 7762
rect 3885 7764 3955 7765
rect 3885 7752 3918 7764
rect 3930 7752 3955 7764
rect 4191 7763 4226 7768
rect 4191 7753 4199 7763
rect 4210 7753 4226 7763
rect 4191 7752 4226 7753
rect 4239 7755 4342 7768
rect 4355 7770 4425 7771
rect 4355 7758 4388 7770
rect 4400 7758 4425 7770
rect 4355 7755 4425 7758
rect 4239 7752 4339 7755
rect 3885 7749 3955 7752
rect 3769 7746 3869 7749
rect 1945 7679 1994 7682
rect 1836 7678 1840 7679
rect 1796 7677 1822 7678
rect 2215 7677 2228 7688
rect 2235 7677 2338 7688
rect 2346 7677 2387 7688
rect 2392 7677 2393 7688
rect 2990 7688 2991 7692
rect 2993 7688 2994 7692
rect 2672 7683 2673 7687
rect 2675 7683 2676 7687
rect 3308 7686 3309 7690
rect 3311 7686 3312 7690
rect 2640 7558 2645 7563
rect 2650 7558 2657 7563
rect 2958 7563 2963 7568
rect 2968 7563 2975 7568
rect 2696 7550 2700 7558
rect 2707 7550 2727 7558
rect 2696 7548 2727 7550
rect 2734 7550 2765 7558
rect 2772 7550 2776 7558
rect 3014 7555 3018 7563
rect 3025 7555 3045 7563
rect 3014 7553 3045 7555
rect 3052 7555 3083 7563
rect 3090 7555 3094 7563
rect 3276 7561 3281 7566
rect 3286 7561 3293 7566
rect 3052 7553 3094 7555
rect 3332 7553 3336 7561
rect 3343 7553 3363 7561
rect 2734 7548 2776 7550
rect 3332 7551 3363 7553
rect 3370 7553 3401 7561
rect 3408 7553 3412 7561
rect 3370 7551 3412 7553
rect 2051 7026 2056 7031
rect 2059 7026 2068 7031
rect 2452 7031 2457 7036
rect 2460 7031 2469 7036
rect 2980 7031 2984 7039
rect 2991 7031 3011 7039
rect 2980 7029 3011 7031
rect 3018 7031 3049 7039
rect 3056 7031 3060 7039
rect 3018 7029 3060 7031
rect 3323 7029 3327 7037
rect 3334 7029 3354 7037
rect 3323 7027 3354 7029
rect 3361 7029 3392 7037
rect 3399 7029 3403 7037
rect 3361 7027 3403 7029
rect 2626 7016 2630 7024
rect 2637 7016 2657 7024
rect 2626 7014 2657 7016
rect 2664 7016 2695 7024
rect 2702 7016 2706 7024
rect 2664 7014 2706 7016
rect 3988 7076 3993 7081
rect 3998 7076 4005 7081
rect 4458 7082 4463 7087
rect 4468 7082 4475 7087
rect 4340 6998 4345 6999
rect 4292 6996 4345 6998
rect 3870 6992 3875 6993
rect 3822 6990 3875 6992
rect 3724 6985 3759 6990
rect 3724 6975 3732 6985
rect 3743 6975 3759 6985
rect 3724 6974 3759 6975
rect 3772 6977 3875 6990
rect 3888 6992 3958 6993
rect 3888 6980 3921 6992
rect 3933 6980 3958 6992
rect 4194 6991 4229 6996
rect 4194 6981 4202 6991
rect 4213 6981 4229 6991
rect 4194 6980 4229 6981
rect 4242 6983 4345 6996
rect 4358 6998 4428 6999
rect 4358 6986 4391 6998
rect 4403 6986 4428 6998
rect 4958 7017 4963 7022
rect 4968 7017 4975 7022
rect 4674 6994 4706 6996
rect 4674 6987 4678 6994
rect 4689 6987 4706 6994
rect 4717 6995 4747 6996
rect 4717 6988 4732 6995
rect 4743 6988 4747 6995
rect 4717 6987 4747 6988
rect 4751 6994 4797 6996
rect 4751 6987 4755 6994
rect 4766 6987 4797 6994
rect 4808 6994 4848 6996
rect 4808 6987 4824 6994
rect 4835 6987 4848 6994
rect 4358 6983 4428 6986
rect 4242 6980 4342 6983
rect 3888 6977 3958 6980
rect 3772 6974 3872 6977
rect 1780 6933 1828 6934
rect 1792 6923 1828 6933
rect 1835 6923 1938 6934
rect 1945 6927 1987 6934
rect 1992 6927 1993 6934
rect 2216 6928 2229 6939
rect 2236 6928 2339 6939
rect 2347 6928 2388 6939
rect 2393 6928 2394 6939
rect 2975 6943 2976 6947
rect 2978 6943 2979 6947
rect 3318 6941 3319 6945
rect 3321 6941 3322 6945
rect 2621 6928 2622 6932
rect 2624 6928 2625 6932
rect 1945 6923 1992 6927
rect 2943 6818 2948 6823
rect 2953 6818 2960 6823
rect 2999 6810 3003 6818
rect 3010 6810 3030 6818
rect 2589 6803 2594 6808
rect 2599 6803 2606 6808
rect 2999 6808 3030 6810
rect 3037 6810 3068 6818
rect 3075 6810 3079 6818
rect 3286 6816 3291 6821
rect 3296 6816 3303 6821
rect 3037 6808 3079 6810
rect 3342 6808 3346 6816
rect 3353 6808 3373 6816
rect 2645 6795 2649 6803
rect 2656 6795 2676 6803
rect 2645 6793 2676 6795
rect 2683 6795 2714 6803
rect 2721 6795 2725 6803
rect 2683 6793 2725 6795
rect 3342 6806 3373 6808
rect 3380 6808 3411 6816
rect 3418 6808 3422 6816
rect 3380 6806 3422 6808
rect 2047 6135 2057 6140
rect 2060 6135 2069 6140
rect 1821 6042 1829 6043
rect 1802 6032 1829 6042
rect 1836 6032 1938 6043
rect 1840 6031 1938 6032
rect 1945 6037 1988 6043
rect 2448 6140 2458 6145
rect 2461 6140 2470 6145
rect 3321 6138 3325 6146
rect 3332 6138 3352 6146
rect 3321 6136 3352 6138
rect 3359 6138 3390 6146
rect 3397 6138 3401 6146
rect 3359 6136 3401 6138
rect 2650 6125 2654 6133
rect 2661 6125 2681 6133
rect 2650 6123 2681 6125
rect 2688 6125 2719 6133
rect 2726 6125 2730 6133
rect 2688 6123 2730 6125
rect 2956 6125 2960 6133
rect 2967 6125 2987 6133
rect 2956 6123 2987 6125
rect 2994 6125 3025 6133
rect 3032 6125 3036 6133
rect 2994 6123 3036 6125
rect 2222 6047 2230 6048
rect 2211 6046 2230 6047
rect 1993 6039 1994 6043
rect 1993 6037 1995 6039
rect 2212 6037 2230 6046
rect 2237 6037 2338 6048
rect 1945 6031 1995 6037
rect 2240 6036 2338 6037
rect 2346 6036 2389 6048
rect 2394 6043 2395 6048
rect 2394 6036 2396 6043
rect 3316 6050 3317 6054
rect 3319 6050 3320 6054
rect 3988 6128 3993 6133
rect 3998 6128 4005 6133
rect 4458 6134 4463 6139
rect 4468 6134 4475 6139
rect 4340 6050 4345 6051
rect 4292 6048 4345 6050
rect 3870 6044 3875 6045
rect 3822 6042 3875 6044
rect 2645 6037 2646 6041
rect 2648 6037 2649 6041
rect 2951 6037 2952 6041
rect 2954 6037 2955 6041
rect 3724 6037 3759 6042
rect 3724 6027 3732 6037
rect 3743 6027 3759 6037
rect 3724 6026 3759 6027
rect 3772 6029 3875 6042
rect 3888 6044 3958 6045
rect 3888 6032 3921 6044
rect 3933 6032 3958 6044
rect 4194 6043 4229 6048
rect 4194 6033 4202 6043
rect 4213 6033 4229 6043
rect 4194 6032 4229 6033
rect 4242 6035 4345 6048
rect 4358 6050 4428 6051
rect 4358 6038 4391 6050
rect 4403 6038 4428 6050
rect 4958 6066 4963 6071
rect 4968 6066 4975 6071
rect 4358 6035 4428 6038
rect 4674 6043 4706 6045
rect 4674 6036 4678 6043
rect 4689 6036 4706 6043
rect 4717 6044 4747 6045
rect 4717 6037 4732 6044
rect 4743 6037 4747 6044
rect 4717 6036 4747 6037
rect 4751 6043 4797 6045
rect 4751 6036 4755 6043
rect 4766 6036 4797 6043
rect 4808 6043 4848 6045
rect 4808 6036 4824 6043
rect 4835 6036 4848 6043
rect 4242 6032 4342 6035
rect 3888 6029 3958 6032
rect 3772 6026 3872 6029
rect 2613 5912 2618 5917
rect 2623 5912 2630 5917
rect 3284 5925 3289 5930
rect 3294 5925 3301 5930
rect 2919 5912 2924 5917
rect 2929 5912 2936 5917
rect 3340 5917 3344 5925
rect 3351 5917 3371 5925
rect 3340 5915 3371 5917
rect 3378 5917 3409 5925
rect 3416 5917 3420 5925
rect 3378 5915 3420 5917
rect 2669 5904 2673 5912
rect 2680 5904 2700 5912
rect 2669 5902 2700 5904
rect 2707 5904 2738 5912
rect 2745 5904 2749 5912
rect 2707 5902 2749 5904
rect 2975 5904 2979 5912
rect 2986 5904 3006 5912
rect 2975 5902 3006 5904
rect 3013 5904 3044 5912
rect 3051 5904 3055 5912
rect 3013 5902 3055 5904
rect 2052 5355 2055 5360
rect 2058 5355 2067 5360
rect 3988 5465 3993 5470
rect 3998 5465 4005 5470
rect 4458 5471 4463 5476
rect 4468 5471 4475 5476
rect 4340 5387 4345 5388
rect 4292 5385 4345 5387
rect 3870 5381 3875 5382
rect 3822 5379 3875 5381
rect 3724 5374 3759 5379
rect 2451 5360 2456 5365
rect 2459 5360 2468 5365
rect 3359 5364 3363 5372
rect 3370 5364 3390 5372
rect 2968 5355 2972 5363
rect 2979 5355 2999 5363
rect 2968 5353 2999 5355
rect 3006 5355 3037 5363
rect 3044 5355 3048 5363
rect 3359 5362 3390 5364
rect 3397 5364 3428 5372
rect 3435 5364 3439 5372
rect 3397 5362 3439 5364
rect 3724 5364 3732 5374
rect 3743 5364 3759 5374
rect 3724 5363 3759 5364
rect 3772 5366 3875 5379
rect 3888 5381 3958 5382
rect 3888 5369 3921 5381
rect 3933 5369 3958 5381
rect 4194 5380 4229 5385
rect 4194 5370 4202 5380
rect 4213 5370 4229 5380
rect 4194 5369 4229 5370
rect 4243 5372 4345 5385
rect 4358 5387 4428 5388
rect 4358 5375 4391 5387
rect 4403 5375 4428 5387
rect 4958 5402 4963 5407
rect 4968 5402 4975 5407
rect 4358 5372 4428 5375
rect 4674 5379 4706 5381
rect 4674 5372 4678 5379
rect 4689 5372 4706 5379
rect 4717 5380 4747 5381
rect 4717 5373 4732 5380
rect 4743 5373 4747 5380
rect 4717 5372 4747 5373
rect 4751 5379 4797 5381
rect 4751 5372 4755 5379
rect 4766 5372 4797 5379
rect 4808 5379 4848 5381
rect 4808 5372 4824 5379
rect 4835 5372 4848 5379
rect 4243 5369 4342 5372
rect 3888 5366 3958 5369
rect 3772 5363 3872 5366
rect 3006 5353 3048 5355
rect 2626 5345 2630 5353
rect 2637 5345 2657 5353
rect 2626 5343 2657 5345
rect 2664 5345 2695 5353
rect 2702 5345 2706 5353
rect 2664 5343 2706 5345
rect 1818 5253 1827 5263
rect 1817 5252 1827 5253
rect 1834 5252 1937 5263
rect 1946 5256 1986 5263
rect 2206 5267 2228 5268
rect 1991 5260 1992 5263
rect 1991 5256 1993 5260
rect 2206 5258 2207 5267
rect 2215 5258 2228 5267
rect 2218 5257 2228 5258
rect 2235 5258 2338 5268
rect 2344 5258 2387 5268
rect 2392 5258 2393 5268
rect 3354 5276 3355 5280
rect 3357 5276 3358 5280
rect 2963 5267 2964 5271
rect 2966 5267 2967 5271
rect 2235 5257 2239 5258
rect 1946 5252 1993 5256
rect 2621 5257 2622 5261
rect 2624 5257 2625 5261
rect 3322 5151 3327 5156
rect 3332 5151 3339 5156
rect 2931 5142 2936 5147
rect 2941 5142 2948 5147
rect 3378 5143 3382 5151
rect 3389 5143 3409 5151
rect 2589 5132 2594 5137
rect 2599 5132 2606 5137
rect 2987 5134 2991 5142
rect 2998 5134 3018 5142
rect 2987 5132 3018 5134
rect 3025 5134 3056 5142
rect 3063 5134 3067 5142
rect 3378 5141 3409 5143
rect 3416 5143 3447 5151
rect 3454 5143 3458 5151
rect 3416 5141 3458 5143
rect 3025 5132 3067 5134
rect 2645 5124 2649 5132
rect 2656 5124 2676 5132
rect 2645 5122 2676 5124
rect 2683 5124 2714 5132
rect 2721 5124 2725 5132
rect 2683 5122 2725 5124
<< pdiffusion >>
rect 1676 8395 1677 8404
rect 1689 8395 1708 8404
rect 1719 8395 1799 8404
rect 1810 8401 1854 8404
rect 1810 8395 1834 8401
rect 1852 8395 1854 8401
rect 1959 8314 1965 8319
rect 1970 8314 1976 8319
rect 1788 7830 1829 7831
rect 1788 7821 1795 7830
rect 1801 7821 1829 7830
rect 1788 7815 1829 7821
rect 1836 7828 1857 7831
rect 1836 7819 1846 7828
rect 1852 7819 1857 7828
rect 1904 7833 1939 7834
rect 1836 7815 1857 7819
rect 1904 7824 1911 7833
rect 1917 7824 1939 7833
rect 1904 7818 1939 7824
rect 1946 7831 1973 7834
rect 1946 7822 1962 7831
rect 1968 7822 1973 7831
rect 2187 7829 2228 7830
rect 1946 7818 1973 7822
rect 2187 7820 2194 7829
rect 2200 7820 2228 7829
rect 2051 7815 2057 7820
rect 2060 7815 2068 7820
rect 2187 7814 2228 7820
rect 2235 7827 2256 7830
rect 2235 7818 2245 7827
rect 2251 7818 2256 7827
rect 2995 7845 3023 7848
rect 2677 7840 2705 7843
rect 2303 7832 2338 7833
rect 2235 7814 2256 7818
rect 2303 7823 2310 7832
rect 2316 7823 2338 7832
rect 2303 7817 2338 7823
rect 2345 7830 2372 7833
rect 2345 7821 2361 7830
rect 2367 7821 2372 7830
rect 2677 7834 2682 7840
rect 2688 7834 2705 7840
rect 2677 7833 2705 7834
rect 2713 7840 2757 7843
rect 2713 7834 2746 7840
rect 2752 7834 2757 7840
rect 2995 7839 3000 7845
rect 3006 7839 3023 7845
rect 2995 7838 3023 7839
rect 3031 7845 3075 7848
rect 3721 7897 3756 7898
rect 3721 7888 3728 7897
rect 3734 7888 3756 7897
rect 3721 7882 3756 7888
rect 3769 7895 3790 7898
rect 3769 7886 3779 7895
rect 3785 7886 3790 7895
rect 3837 7900 3872 7901
rect 3769 7882 3790 7886
rect 3837 7891 3844 7900
rect 3850 7891 3872 7900
rect 3837 7885 3872 7891
rect 3889 7898 3906 7901
rect 3889 7889 3895 7898
rect 3901 7889 3906 7898
rect 4191 7903 4226 7904
rect 4191 7894 4198 7903
rect 4204 7894 4226 7903
rect 3889 7885 3906 7889
rect 4191 7888 4226 7894
rect 4239 7901 4260 7904
rect 4239 7892 4249 7901
rect 4255 7892 4260 7901
rect 4674 7934 4675 7943
rect 4687 7934 4706 7943
rect 4717 7934 4797 7943
rect 4808 7940 4852 7943
rect 4808 7934 4832 7940
rect 4850 7934 4852 7940
rect 4307 7906 4341 7907
rect 4239 7888 4260 7892
rect 4307 7897 4314 7906
rect 4320 7897 4341 7906
rect 4307 7891 4341 7897
rect 4357 7904 4376 7907
rect 4357 7895 4365 7904
rect 4371 7895 4376 7904
rect 4357 7891 4376 7895
rect 3031 7839 3064 7845
rect 3070 7839 3075 7845
rect 3031 7838 3075 7839
rect 3313 7843 3341 7846
rect 3313 7837 3318 7843
rect 3324 7837 3341 7843
rect 3313 7836 3341 7837
rect 3349 7843 3393 7846
rect 3349 7837 3382 7843
rect 3388 7837 3393 7843
rect 3349 7836 3393 7837
rect 2713 7833 2757 7834
rect 2345 7817 2372 7821
rect 2450 7814 2456 7819
rect 2459 7814 2467 7819
rect 3984 7882 3990 7887
rect 3995 7882 4001 7887
rect 4454 7888 4460 7893
rect 4465 7888 4471 7893
rect 4957 7853 4963 7858
rect 4968 7853 4974 7858
rect 2990 7708 2991 7712
rect 2993 7708 2994 7712
rect 2672 7703 2673 7707
rect 2675 7703 2676 7707
rect 3308 7706 3309 7710
rect 3311 7706 3312 7710
rect 1787 7075 1828 7076
rect 1787 7066 1794 7075
rect 1800 7066 1828 7075
rect 1787 7060 1828 7066
rect 1835 7073 1856 7076
rect 1835 7064 1845 7073
rect 1851 7064 1856 7073
rect 1903 7078 1938 7079
rect 1835 7060 1856 7064
rect 1903 7069 1910 7078
rect 1916 7069 1938 7078
rect 1903 7063 1938 7069
rect 1945 7076 1972 7079
rect 1945 7067 1961 7076
rect 1967 7067 1972 7076
rect 2188 7080 2229 7081
rect 1945 7063 1972 7067
rect 2188 7071 2195 7080
rect 2201 7071 2229 7080
rect 2188 7065 2229 7071
rect 2236 7078 2257 7081
rect 2236 7069 2246 7078
rect 2252 7069 2257 7078
rect 3014 7624 3041 7627
rect 2696 7619 2723 7622
rect 2696 7613 2701 7619
rect 2707 7613 2723 7619
rect 2696 7612 2723 7613
rect 2736 7619 2776 7622
rect 2736 7613 2765 7619
rect 2771 7613 2776 7619
rect 3014 7618 3019 7624
rect 3025 7618 3041 7624
rect 3014 7617 3041 7618
rect 3054 7624 3094 7627
rect 3054 7618 3083 7624
rect 3089 7618 3094 7624
rect 3054 7617 3094 7618
rect 3332 7622 3359 7625
rect 3332 7616 3337 7622
rect 3343 7616 3359 7622
rect 3332 7615 3359 7616
rect 3372 7622 3412 7625
rect 3372 7616 3401 7622
rect 3407 7616 3412 7622
rect 3372 7615 3412 7616
rect 2736 7612 2776 7613
rect 2957 7597 2963 7602
rect 2968 7597 2974 7602
rect 2639 7592 2645 7597
rect 2650 7592 2656 7597
rect 3275 7595 3281 7600
rect 3286 7595 3292 7600
rect 2304 7083 2339 7084
rect 2236 7065 2257 7069
rect 2304 7074 2311 7083
rect 2317 7074 2339 7083
rect 2304 7068 2339 7074
rect 2346 7081 2373 7084
rect 2346 7072 2362 7081
rect 2368 7072 2373 7081
rect 2980 7100 3008 7103
rect 2980 7094 2985 7100
rect 2991 7094 3008 7100
rect 2980 7093 3008 7094
rect 3016 7100 3060 7103
rect 3724 7125 3758 7126
rect 3724 7116 3731 7125
rect 3737 7116 3758 7125
rect 3724 7110 3758 7116
rect 3772 7123 3793 7126
rect 3772 7114 3782 7123
rect 3788 7114 3793 7123
rect 3840 7128 3875 7129
rect 3772 7110 3793 7114
rect 3840 7119 3847 7128
rect 3853 7119 3875 7128
rect 3840 7113 3875 7119
rect 3888 7126 3909 7129
rect 3888 7117 3898 7126
rect 3904 7117 3909 7126
rect 4194 7131 4229 7132
rect 4194 7122 4201 7131
rect 4207 7122 4229 7131
rect 3888 7113 3909 7117
rect 4194 7116 4229 7122
rect 4242 7129 4263 7132
rect 4242 7120 4252 7129
rect 4258 7120 4263 7129
rect 4310 7134 4345 7135
rect 4242 7116 4263 7120
rect 4310 7125 4317 7134
rect 4323 7125 4345 7134
rect 4310 7119 4345 7125
rect 4358 7132 4379 7135
rect 4358 7123 4368 7132
rect 4374 7123 4379 7132
rect 4674 7132 4675 7141
rect 4687 7132 4706 7141
rect 4717 7132 4797 7141
rect 4808 7138 4852 7141
rect 4808 7132 4832 7138
rect 4850 7132 4852 7138
rect 4358 7119 4379 7123
rect 3016 7094 3049 7100
rect 3055 7094 3060 7100
rect 3016 7093 3060 7094
rect 3323 7098 3351 7101
rect 3323 7092 3328 7098
rect 3334 7092 3351 7098
rect 3323 7091 3351 7092
rect 3359 7098 3403 7101
rect 3359 7092 3392 7098
rect 3398 7092 3403 7098
rect 3359 7091 3403 7092
rect 2626 7085 2654 7088
rect 2626 7079 2631 7085
rect 2637 7079 2654 7085
rect 2626 7078 2654 7079
rect 2662 7085 2706 7088
rect 2662 7079 2695 7085
rect 2701 7079 2706 7085
rect 2662 7078 2706 7079
rect 2346 7068 2373 7072
rect 2050 7060 2056 7065
rect 2059 7060 2067 7065
rect 2451 7065 2457 7070
rect 2460 7065 2468 7070
rect 3987 7110 3993 7115
rect 3998 7110 4004 7115
rect 4457 7116 4463 7121
rect 4468 7116 4474 7121
rect 4957 7051 4963 7056
rect 4968 7051 4974 7056
rect 2975 6963 2976 6967
rect 2978 6963 2979 6967
rect 2621 6948 2622 6952
rect 2624 6948 2625 6952
rect 3318 6961 3319 6965
rect 3321 6961 3322 6965
rect 1788 6184 1829 6185
rect 1788 6175 1795 6184
rect 1801 6175 1829 6184
rect 1788 6169 1829 6175
rect 1836 6182 1857 6185
rect 1836 6173 1846 6182
rect 1852 6173 1857 6182
rect 1904 6187 1938 6188
rect 1836 6169 1857 6173
rect 1904 6178 1911 6187
rect 1917 6178 1938 6187
rect 1904 6172 1938 6178
rect 1945 6185 1973 6188
rect 1945 6176 1962 6185
rect 1968 6176 1973 6185
rect 2189 6189 2230 6190
rect 1945 6172 1973 6176
rect 2189 6180 2196 6189
rect 2202 6180 2230 6189
rect 2189 6174 2230 6180
rect 2237 6187 2258 6190
rect 2237 6178 2247 6187
rect 2253 6178 2258 6187
rect 2999 6879 3026 6882
rect 2999 6873 3004 6879
rect 3010 6873 3026 6879
rect 2999 6872 3026 6873
rect 3039 6879 3079 6882
rect 3039 6873 3068 6879
rect 3074 6873 3079 6879
rect 3039 6872 3079 6873
rect 3342 6877 3369 6880
rect 3342 6871 3347 6877
rect 3353 6871 3369 6877
rect 3342 6870 3369 6871
rect 3382 6877 3422 6880
rect 3382 6871 3411 6877
rect 3417 6871 3422 6877
rect 3382 6870 3422 6871
rect 2645 6864 2672 6867
rect 2645 6858 2650 6864
rect 2656 6858 2672 6864
rect 2645 6857 2672 6858
rect 2685 6864 2725 6867
rect 2685 6858 2714 6864
rect 2720 6858 2725 6864
rect 2685 6857 2725 6858
rect 2942 6852 2948 6857
rect 2953 6852 2959 6857
rect 2588 6837 2594 6842
rect 2599 6837 2605 6842
rect 3285 6850 3291 6855
rect 3296 6850 3302 6855
rect 2305 6192 2340 6193
rect 2237 6174 2258 6178
rect 2305 6183 2312 6192
rect 2318 6183 2340 6192
rect 2305 6177 2340 6183
rect 2347 6190 2374 6193
rect 2347 6181 2363 6190
rect 2369 6181 2374 6190
rect 3321 6207 3349 6210
rect 3321 6201 3326 6207
rect 3332 6201 3349 6207
rect 3321 6200 3349 6201
rect 3357 6207 3401 6210
rect 3357 6201 3390 6207
rect 3396 6201 3401 6207
rect 3357 6200 3401 6201
rect 2650 6194 2678 6197
rect 2650 6188 2655 6194
rect 2661 6188 2678 6194
rect 2650 6187 2678 6188
rect 2686 6194 2730 6197
rect 2686 6188 2719 6194
rect 2725 6188 2730 6194
rect 2686 6187 2730 6188
rect 2956 6194 2984 6197
rect 2956 6188 2961 6194
rect 2967 6188 2984 6194
rect 2956 6187 2984 6188
rect 2992 6194 3036 6197
rect 2992 6188 3025 6194
rect 3031 6188 3036 6194
rect 2992 6187 3036 6188
rect 2347 6177 2374 6181
rect 2051 6169 2057 6174
rect 2060 6169 2068 6174
rect 2452 6174 2458 6179
rect 2461 6174 2469 6179
rect 3724 6177 3759 6178
rect 3724 6168 3731 6177
rect 3737 6168 3759 6177
rect 3724 6162 3759 6168
rect 3772 6175 3793 6178
rect 3772 6166 3782 6175
rect 3788 6166 3793 6175
rect 3840 6180 3875 6181
rect 3772 6162 3793 6166
rect 3840 6171 3847 6180
rect 3853 6171 3875 6180
rect 3840 6165 3875 6171
rect 3891 6178 3909 6181
rect 3891 6169 3898 6178
rect 3904 6169 3909 6178
rect 4194 6183 4229 6184
rect 4194 6174 4201 6183
rect 4207 6174 4229 6183
rect 3891 6165 3909 6169
rect 4194 6168 4229 6174
rect 4242 6181 4263 6184
rect 4242 6172 4252 6181
rect 4258 6172 4263 6181
rect 4310 6186 4344 6187
rect 4242 6168 4263 6172
rect 4310 6177 4317 6186
rect 4323 6177 4344 6186
rect 4310 6171 4344 6177
rect 4360 6184 4379 6187
rect 4360 6175 4368 6184
rect 4374 6175 4379 6184
rect 4674 6181 4675 6190
rect 4687 6181 4706 6190
rect 4717 6181 4797 6190
rect 4808 6187 4852 6190
rect 4808 6181 4832 6187
rect 4850 6181 4852 6187
rect 4360 6171 4379 6175
rect 3316 6070 3317 6074
rect 3319 6070 3320 6074
rect 2645 6057 2646 6061
rect 2648 6057 2649 6061
rect 2951 6057 2952 6061
rect 2954 6057 2955 6061
rect 1786 5404 1827 5405
rect 1786 5395 1793 5404
rect 1799 5395 1827 5404
rect 1786 5389 1827 5395
rect 1834 5402 1855 5405
rect 1834 5393 1844 5402
rect 1850 5393 1855 5402
rect 3987 6162 3993 6167
rect 3998 6162 4004 6167
rect 4457 6168 4463 6173
rect 4468 6168 4474 6173
rect 1902 5407 1937 5408
rect 1834 5389 1855 5393
rect 1902 5398 1909 5407
rect 1915 5398 1937 5407
rect 1902 5392 1937 5398
rect 1945 5405 1971 5408
rect 1945 5396 1960 5405
rect 1966 5396 1971 5405
rect 2187 5409 2228 5410
rect 1945 5392 1971 5396
rect 2187 5400 2194 5409
rect 2200 5400 2228 5409
rect 2187 5394 2228 5400
rect 2235 5407 2256 5410
rect 2235 5398 2245 5407
rect 2251 5398 2256 5407
rect 4957 6100 4963 6105
rect 4968 6100 4974 6105
rect 3340 5986 3367 5989
rect 3340 5980 3345 5986
rect 3351 5980 3367 5986
rect 3340 5979 3367 5980
rect 3380 5986 3420 5989
rect 3380 5980 3409 5986
rect 3415 5980 3420 5986
rect 3380 5979 3420 5980
rect 2669 5973 2696 5976
rect 2669 5967 2674 5973
rect 2680 5967 2696 5973
rect 2669 5966 2696 5967
rect 2709 5973 2749 5976
rect 2709 5967 2738 5973
rect 2744 5967 2749 5973
rect 2709 5966 2749 5967
rect 2975 5973 3002 5976
rect 2975 5967 2980 5973
rect 2986 5967 3002 5973
rect 2975 5966 3002 5967
rect 3015 5973 3055 5976
rect 3015 5967 3044 5973
rect 3050 5967 3055 5973
rect 3015 5966 3055 5967
rect 3283 5959 3289 5964
rect 3294 5959 3300 5964
rect 2612 5946 2618 5951
rect 2623 5946 2629 5951
rect 2918 5946 2924 5951
rect 2929 5946 2935 5951
rect 3724 5514 3759 5515
rect 3724 5505 3731 5514
rect 3737 5505 3759 5514
rect 3724 5499 3759 5505
rect 3772 5512 3793 5515
rect 3772 5503 3782 5512
rect 3788 5503 3793 5512
rect 3840 5517 3873 5518
rect 3772 5499 3793 5503
rect 3840 5508 3847 5517
rect 3853 5508 3873 5517
rect 3840 5502 3873 5508
rect 3888 5515 3909 5518
rect 3888 5506 3898 5515
rect 3904 5506 3909 5515
rect 4194 5520 4229 5521
rect 4194 5511 4201 5520
rect 4207 5511 4229 5520
rect 3888 5502 3909 5506
rect 4194 5505 4229 5511
rect 4242 5518 4263 5521
rect 4242 5509 4252 5518
rect 4258 5509 4263 5518
rect 4310 5523 4345 5524
rect 4242 5505 4263 5509
rect 4310 5514 4317 5523
rect 4323 5514 4345 5523
rect 4310 5508 4345 5514
rect 4361 5521 4379 5524
rect 4361 5512 4368 5521
rect 4374 5512 4379 5521
rect 4674 5517 4675 5526
rect 4687 5517 4706 5526
rect 4717 5517 4797 5526
rect 4808 5523 4852 5526
rect 4808 5517 4832 5523
rect 4850 5517 4852 5523
rect 4361 5508 4379 5512
rect 2303 5412 2338 5413
rect 2235 5394 2256 5398
rect 2303 5403 2310 5412
rect 2316 5403 2338 5412
rect 2303 5397 2338 5403
rect 2345 5410 2372 5413
rect 2345 5401 2361 5410
rect 2367 5401 2372 5410
rect 3359 5433 3387 5436
rect 3359 5427 3364 5433
rect 3370 5427 3387 5433
rect 2968 5424 2996 5427
rect 2968 5418 2973 5424
rect 2979 5418 2996 5424
rect 2968 5417 2996 5418
rect 3004 5424 3048 5427
rect 3359 5426 3387 5427
rect 3395 5433 3439 5436
rect 3395 5427 3428 5433
rect 3434 5427 3439 5433
rect 3395 5426 3439 5427
rect 3004 5418 3037 5424
rect 3043 5418 3048 5424
rect 3004 5417 3048 5418
rect 2626 5414 2654 5417
rect 2626 5408 2631 5414
rect 2637 5408 2654 5414
rect 2626 5407 2654 5408
rect 2662 5414 2706 5417
rect 2662 5408 2695 5414
rect 2701 5408 2706 5414
rect 2662 5407 2706 5408
rect 2345 5397 2372 5401
rect 2049 5389 2055 5394
rect 2058 5389 2066 5394
rect 2450 5394 2456 5399
rect 2459 5394 2467 5399
rect 3987 5499 3993 5504
rect 3998 5499 4004 5504
rect 4457 5505 4463 5510
rect 4468 5505 4474 5510
rect 4957 5436 4963 5441
rect 4968 5436 4974 5441
rect 3354 5296 3355 5300
rect 3357 5296 3358 5300
rect 2963 5287 2964 5291
rect 2966 5287 2967 5291
rect 2621 5277 2622 5281
rect 2624 5277 2625 5281
rect 3378 5212 3405 5215
rect 3378 5206 3383 5212
rect 3389 5206 3405 5212
rect 2987 5203 3014 5206
rect 2987 5197 2992 5203
rect 2998 5197 3014 5203
rect 2987 5196 3014 5197
rect 3027 5203 3067 5206
rect 3378 5205 3405 5206
rect 3418 5212 3458 5215
rect 3418 5206 3447 5212
rect 3453 5206 3458 5212
rect 3418 5205 3458 5206
rect 3027 5197 3056 5203
rect 3062 5197 3067 5203
rect 3027 5196 3067 5197
rect 2645 5193 2672 5196
rect 2645 5187 2650 5193
rect 2656 5187 2672 5193
rect 2645 5186 2672 5187
rect 2685 5193 2725 5196
rect 2685 5187 2714 5193
rect 2720 5187 2725 5193
rect 2685 5186 2725 5187
rect 3321 5185 3327 5190
rect 3332 5185 3338 5190
rect 2930 5176 2936 5181
rect 2941 5176 2947 5181
rect 2588 5166 2594 5171
rect 2599 5166 2605 5171
<< ndcontact >>
rect 1954 8280 1960 8285
rect 1977 8280 1983 8285
rect 1680 8250 1691 8257
rect 1734 8251 1745 8258
rect 1757 8250 1768 8257
rect 1826 8250 1837 8257
rect 2043 7781 2051 7786
rect 2069 7781 2075 7786
rect 1769 7677 1796 7688
rect 1988 7682 1993 7694
rect 2443 7779 2451 7785
rect 2468 7780 2474 7785
rect 2681 7771 2688 7779
rect 2746 7771 2753 7779
rect 2999 7776 3006 7784
rect 3064 7776 3071 7784
rect 3317 7774 3324 7782
rect 3382 7774 3389 7782
rect 3979 7848 3985 7853
rect 4002 7848 4008 7853
rect 4449 7854 4455 7859
rect 4472 7854 4478 7859
rect 4952 7819 4958 7824
rect 4975 7819 4981 7824
rect 4678 7789 4689 7796
rect 4732 7790 4743 7797
rect 4755 7789 4766 7796
rect 4824 7789 4835 7796
rect 3729 7747 3740 7757
rect 3918 7752 3930 7764
rect 4199 7753 4210 7763
rect 4388 7758 4400 7770
rect 2197 7676 2215 7688
rect 2387 7677 2392 7688
rect 2986 7688 2990 7692
rect 2994 7688 2998 7692
rect 2668 7683 2672 7687
rect 2676 7683 2680 7687
rect 3304 7686 3308 7690
rect 3312 7686 3316 7690
rect 2634 7558 2640 7563
rect 2657 7558 2663 7563
rect 2952 7563 2958 7568
rect 2975 7563 2981 7568
rect 2700 7550 2707 7558
rect 2765 7550 2772 7558
rect 3018 7555 3025 7563
rect 3083 7555 3090 7563
rect 3270 7561 3276 7566
rect 3293 7561 3299 7566
rect 3336 7553 3343 7561
rect 3401 7553 3408 7561
rect 2044 7025 2051 7031
rect 2068 7026 2074 7031
rect 2444 7030 2452 7036
rect 2469 7031 2475 7036
rect 2984 7031 2991 7039
rect 3049 7031 3056 7039
rect 3327 7029 3334 7037
rect 3392 7029 3399 7037
rect 2630 7016 2637 7024
rect 2695 7016 2702 7024
rect 3982 7076 3988 7081
rect 4005 7076 4011 7081
rect 4452 7082 4458 7087
rect 4475 7082 4481 7087
rect 3732 6975 3743 6985
rect 3921 6980 3933 6992
rect 4202 6981 4213 6991
rect 4391 6986 4403 6998
rect 4952 7017 4958 7022
rect 4975 7017 4981 7022
rect 4678 6987 4689 6994
rect 4732 6988 4743 6995
rect 4755 6987 4766 6994
rect 4824 6987 4835 6994
rect 1779 6923 1792 6933
rect 1987 6927 1992 6939
rect 2198 6927 2216 6939
rect 2388 6928 2393 6939
rect 2971 6943 2975 6947
rect 2979 6943 2983 6947
rect 3314 6941 3318 6945
rect 3322 6941 3326 6945
rect 2617 6928 2621 6932
rect 2625 6928 2629 6932
rect 2937 6818 2943 6823
rect 2960 6818 2966 6823
rect 3003 6810 3010 6818
rect 2583 6803 2589 6808
rect 2606 6803 2612 6808
rect 3068 6810 3075 6818
rect 3280 6816 3286 6821
rect 3303 6816 3309 6821
rect 3346 6808 3353 6816
rect 2649 6795 2656 6803
rect 2714 6795 2721 6803
rect 3411 6808 3418 6816
rect 2043 6135 2047 6140
rect 2069 6135 2075 6140
rect 1787 6031 1802 6042
rect 1988 6037 1993 6049
rect 2444 6139 2448 6145
rect 2470 6140 2476 6145
rect 3325 6138 3332 6146
rect 3390 6138 3397 6146
rect 2654 6125 2661 6133
rect 2719 6125 2726 6133
rect 2960 6125 2967 6133
rect 3025 6125 3032 6133
rect 2202 6037 2212 6046
rect 2389 6035 2394 6048
rect 3312 6050 3316 6054
rect 3320 6050 3324 6054
rect 3982 6128 3988 6133
rect 4005 6128 4011 6133
rect 4452 6134 4458 6139
rect 4475 6134 4481 6139
rect 2641 6037 2645 6041
rect 2649 6037 2653 6041
rect 2947 6037 2951 6041
rect 2955 6037 2959 6041
rect 3732 6027 3743 6037
rect 3921 6032 3933 6044
rect 4202 6033 4213 6043
rect 4391 6038 4403 6050
rect 4952 6066 4958 6071
rect 4975 6066 4981 6071
rect 4678 6036 4689 6043
rect 4732 6037 4743 6044
rect 4755 6036 4766 6043
rect 4824 6036 4835 6043
rect 2607 5912 2613 5917
rect 2630 5912 2636 5917
rect 3278 5925 3284 5930
rect 3301 5925 3307 5930
rect 2913 5912 2919 5917
rect 2936 5912 2942 5917
rect 3344 5917 3351 5925
rect 3409 5917 3416 5925
rect 2673 5904 2680 5912
rect 2738 5904 2745 5912
rect 2979 5904 2986 5912
rect 3044 5904 3051 5912
rect 2044 5355 2052 5360
rect 2067 5355 2073 5360
rect 3982 5465 3988 5470
rect 4005 5465 4011 5470
rect 4452 5471 4458 5476
rect 4475 5471 4481 5476
rect 2444 5359 2451 5365
rect 2468 5360 2474 5365
rect 3363 5364 3370 5372
rect 2972 5355 2979 5363
rect 3037 5355 3044 5363
rect 3428 5364 3435 5372
rect 3732 5364 3743 5374
rect 3921 5369 3933 5381
rect 4202 5370 4213 5380
rect 4391 5375 4403 5387
rect 4952 5402 4958 5407
rect 4975 5402 4981 5407
rect 4678 5372 4689 5379
rect 4732 5373 4743 5380
rect 4755 5372 4766 5379
rect 4824 5372 4835 5379
rect 2630 5345 2637 5353
rect 2695 5345 2702 5353
rect 1804 5253 1818 5263
rect 1986 5256 1991 5268
rect 2207 5258 2215 5267
rect 2387 5258 2392 5268
rect 3350 5276 3354 5280
rect 3358 5276 3362 5280
rect 2959 5267 2963 5271
rect 2967 5267 2971 5271
rect 2617 5257 2621 5261
rect 2625 5257 2629 5261
rect 3316 5151 3322 5156
rect 3339 5151 3345 5156
rect 2925 5142 2931 5147
rect 2948 5142 2954 5147
rect 3382 5143 3389 5151
rect 2583 5132 2589 5137
rect 2606 5132 2612 5137
rect 2991 5134 2998 5142
rect 3056 5134 3063 5142
rect 3447 5143 3454 5151
rect 2649 5124 2656 5132
rect 2714 5124 2721 5132
<< pdcontact >>
rect 1677 8395 1689 8404
rect 1834 8395 1852 8401
rect 1953 8314 1959 8319
rect 1976 8314 1982 8319
rect 1795 7821 1801 7830
rect 1846 7819 1852 7828
rect 1911 7824 1917 7833
rect 1962 7822 1968 7831
rect 2194 7820 2200 7829
rect 2045 7815 2051 7820
rect 2068 7815 2074 7820
rect 2245 7818 2251 7827
rect 2310 7823 2316 7832
rect 2361 7821 2367 7830
rect 2682 7834 2688 7840
rect 2746 7834 2752 7840
rect 3000 7839 3006 7845
rect 3728 7888 3734 7897
rect 3779 7886 3785 7895
rect 3844 7891 3850 7900
rect 3895 7889 3901 7898
rect 4198 7894 4204 7903
rect 4249 7892 4255 7901
rect 4675 7934 4687 7943
rect 4832 7934 4850 7940
rect 4314 7897 4320 7906
rect 4365 7895 4371 7904
rect 3064 7839 3070 7845
rect 3318 7837 3324 7843
rect 3382 7837 3388 7843
rect 2444 7814 2450 7819
rect 2467 7814 2473 7819
rect 3978 7882 3984 7887
rect 4001 7882 4007 7887
rect 4448 7888 4454 7893
rect 4471 7888 4477 7893
rect 4951 7853 4957 7858
rect 4974 7853 4980 7858
rect 2986 7708 2990 7712
rect 2994 7708 2998 7712
rect 2668 7703 2672 7707
rect 2676 7703 2680 7707
rect 3304 7706 3308 7710
rect 3312 7706 3316 7710
rect 1794 7066 1800 7075
rect 1845 7064 1851 7073
rect 1910 7069 1916 7078
rect 1961 7067 1967 7076
rect 2195 7071 2201 7080
rect 2246 7069 2252 7078
rect 2701 7613 2707 7619
rect 2765 7613 2771 7619
rect 3019 7618 3025 7624
rect 3083 7618 3089 7624
rect 3337 7616 3343 7622
rect 3401 7616 3407 7622
rect 2951 7597 2957 7602
rect 2974 7597 2980 7602
rect 2633 7592 2639 7597
rect 2656 7592 2662 7597
rect 3269 7595 3275 7600
rect 3292 7595 3298 7600
rect 2311 7074 2317 7083
rect 2362 7072 2368 7081
rect 2985 7094 2991 7100
rect 3731 7116 3737 7125
rect 3782 7114 3788 7123
rect 3847 7119 3853 7128
rect 3898 7117 3904 7126
rect 4201 7122 4207 7131
rect 4252 7120 4258 7129
rect 4317 7125 4323 7134
rect 4368 7123 4374 7132
rect 4675 7132 4687 7141
rect 4832 7132 4850 7138
rect 3049 7094 3055 7100
rect 3328 7092 3334 7098
rect 3392 7092 3398 7098
rect 2631 7079 2637 7085
rect 2695 7079 2701 7085
rect 2044 7060 2050 7065
rect 2067 7060 2073 7065
rect 2445 7065 2451 7070
rect 2468 7065 2474 7070
rect 3981 7110 3987 7115
rect 4004 7110 4010 7115
rect 4451 7116 4457 7121
rect 4474 7116 4480 7121
rect 4951 7051 4957 7056
rect 4974 7051 4980 7056
rect 2971 6963 2975 6967
rect 2979 6963 2983 6967
rect 2617 6948 2621 6952
rect 2625 6948 2629 6952
rect 3314 6961 3318 6965
rect 3322 6961 3326 6965
rect 1795 6175 1801 6184
rect 1846 6173 1852 6182
rect 1911 6178 1917 6187
rect 1962 6176 1968 6185
rect 2196 6180 2202 6189
rect 2247 6178 2253 6187
rect 3004 6873 3010 6879
rect 3068 6873 3074 6879
rect 3347 6871 3353 6877
rect 3411 6871 3417 6877
rect 2650 6858 2656 6864
rect 2714 6858 2720 6864
rect 2936 6852 2942 6857
rect 2959 6852 2965 6857
rect 2582 6837 2588 6842
rect 2605 6837 2611 6842
rect 3279 6850 3285 6855
rect 3302 6850 3308 6855
rect 2312 6183 2318 6192
rect 2363 6181 2369 6190
rect 3326 6201 3332 6207
rect 3390 6201 3396 6207
rect 2655 6188 2661 6194
rect 2719 6188 2725 6194
rect 2961 6188 2967 6194
rect 3025 6188 3031 6194
rect 2045 6169 2051 6174
rect 2068 6169 2074 6174
rect 2446 6174 2452 6179
rect 2469 6174 2475 6179
rect 3731 6168 3737 6177
rect 3782 6166 3788 6175
rect 3847 6171 3853 6180
rect 3898 6169 3904 6178
rect 4201 6174 4207 6183
rect 4252 6172 4258 6181
rect 4317 6177 4323 6186
rect 4368 6175 4374 6184
rect 4675 6181 4687 6190
rect 4832 6181 4850 6187
rect 3312 6070 3316 6074
rect 3320 6070 3324 6074
rect 2641 6057 2645 6061
rect 2649 6057 2653 6061
rect 2947 6057 2951 6061
rect 2955 6057 2959 6061
rect 1793 5395 1799 5404
rect 1844 5393 1850 5402
rect 3981 6162 3987 6167
rect 4004 6162 4010 6167
rect 4451 6168 4457 6173
rect 4474 6168 4480 6173
rect 1909 5398 1915 5407
rect 1960 5396 1966 5405
rect 2194 5400 2200 5409
rect 2245 5398 2251 5407
rect 4951 6100 4957 6105
rect 4974 6100 4980 6105
rect 3345 5980 3351 5986
rect 3409 5980 3415 5986
rect 2674 5967 2680 5973
rect 2738 5967 2744 5973
rect 2980 5967 2986 5973
rect 3044 5967 3050 5973
rect 3277 5959 3283 5964
rect 3300 5959 3306 5964
rect 2606 5946 2612 5951
rect 2629 5946 2635 5951
rect 2912 5946 2918 5951
rect 2935 5946 2941 5951
rect 3731 5505 3737 5514
rect 3782 5503 3788 5512
rect 3847 5508 3853 5517
rect 3898 5506 3904 5515
rect 4201 5511 4207 5520
rect 4252 5509 4258 5518
rect 4317 5514 4323 5523
rect 4368 5512 4374 5521
rect 4675 5517 4687 5526
rect 4832 5517 4850 5523
rect 2310 5403 2316 5412
rect 2361 5401 2367 5410
rect 3364 5427 3370 5433
rect 2973 5418 2979 5424
rect 3428 5427 3434 5433
rect 3037 5418 3043 5424
rect 2631 5408 2637 5414
rect 2695 5408 2701 5414
rect 2043 5389 2049 5394
rect 2066 5389 2072 5394
rect 2444 5394 2450 5399
rect 2467 5394 2473 5399
rect 3981 5499 3987 5504
rect 4004 5499 4010 5504
rect 4451 5505 4457 5510
rect 4474 5505 4480 5510
rect 4951 5436 4957 5441
rect 4974 5436 4980 5441
rect 3350 5296 3354 5300
rect 3358 5296 3362 5300
rect 2959 5287 2963 5291
rect 2967 5287 2971 5291
rect 2617 5277 2621 5281
rect 2625 5277 2629 5281
rect 3383 5206 3389 5212
rect 2992 5197 2998 5203
rect 3447 5206 3453 5212
rect 3056 5197 3062 5203
rect 2650 5187 2656 5193
rect 2714 5187 2720 5193
rect 3315 5185 3321 5190
rect 3338 5185 3344 5190
rect 2924 5176 2930 5181
rect 2947 5176 2953 5181
rect 2582 5166 2588 5171
rect 2605 5166 2611 5171
<< nsubstratencontact >>
rect 1869 8389 1881 8405
rect 1941 8319 1945 8326
rect 1870 7825 1881 7843
rect 1985 7823 1996 7841
rect 2033 7820 2037 7827
rect 2269 7824 2280 7842
rect 2674 7863 2689 7874
rect 2992 7868 3007 7879
rect 3310 7866 3325 7877
rect 2384 7822 2395 7840
rect 3803 7892 3814 7910
rect 3918 7890 3929 7908
rect 3966 7887 3970 7894
rect 4273 7898 4284 7916
rect 4388 7896 4399 7914
rect 4436 7893 4440 7900
rect 2432 7819 2436 7826
rect 4867 7928 4879 7944
rect 4939 7858 4943 7865
rect 2686 7709 2692 7715
rect 3004 7714 3010 7720
rect 3322 7712 3328 7718
rect 1869 7070 1880 7088
rect 1984 7068 1995 7086
rect 2032 7065 2036 7072
rect 2270 7075 2281 7093
rect 2687 7641 2702 7649
rect 3005 7646 3020 7654
rect 3323 7644 3338 7652
rect 2621 7597 2625 7604
rect 2939 7602 2943 7609
rect 3257 7600 3261 7607
rect 2623 7108 2638 7119
rect 2385 7073 2396 7091
rect 2977 7123 2992 7134
rect 3320 7121 3335 7132
rect 3806 7120 3817 7138
rect 3921 7118 3932 7136
rect 3969 7115 3973 7122
rect 4276 7126 4287 7144
rect 4391 7124 4402 7142
rect 4439 7121 4443 7128
rect 2433 7070 2437 7077
rect 4867 7126 4879 7142
rect 4939 7056 4943 7063
rect 2989 6969 2995 6975
rect 3332 6967 3338 6973
rect 2635 6954 2641 6960
rect 1870 6179 1881 6197
rect 1985 6177 1996 6195
rect 2033 6174 2037 6181
rect 2271 6184 2282 6202
rect 2636 6886 2651 6894
rect 2990 6901 3005 6909
rect 3333 6899 3348 6907
rect 2924 6857 2928 6864
rect 3267 6855 3271 6862
rect 2570 6842 2574 6849
rect 2647 6217 2662 6228
rect 2386 6182 2397 6200
rect 2953 6217 2968 6228
rect 3318 6230 3333 6241
rect 2434 6179 2438 6186
rect 3806 6172 3817 6190
rect 3921 6170 3932 6188
rect 3969 6167 3973 6174
rect 4276 6178 4287 6196
rect 4391 6176 4402 6194
rect 4439 6173 4443 6180
rect 3330 6076 3336 6082
rect 2659 6063 2665 6069
rect 2965 6063 2971 6069
rect 1868 5399 1879 5417
rect 4867 6175 4879 6191
rect 1983 5397 1994 5415
rect 2031 5394 2035 5401
rect 2269 5404 2280 5422
rect 4939 6105 4943 6112
rect 2660 5995 2675 6003
rect 2966 5995 2981 6003
rect 3331 6008 3346 6016
rect 3265 5964 3269 5971
rect 2594 5951 2598 5958
rect 2900 5951 2904 5958
rect 3806 5509 3817 5527
rect 3921 5507 3932 5525
rect 3969 5504 3973 5511
rect 4276 5515 4287 5533
rect 4391 5513 4402 5531
rect 4439 5510 4443 5517
rect 2623 5437 2638 5448
rect 2384 5402 2395 5420
rect 2965 5447 2980 5458
rect 3356 5456 3371 5467
rect 2432 5399 2436 5406
rect 4867 5511 4879 5527
rect 4939 5441 4943 5448
rect 3368 5302 3374 5308
rect 2977 5293 2983 5299
rect 2635 5283 2641 5289
rect 2636 5215 2651 5223
rect 2978 5225 2993 5233
rect 3369 5234 3384 5242
rect 3303 5190 3307 5197
rect 2912 5181 2916 5188
rect 2570 5171 2574 5178
<< polysilicon >>
rect 1708 8404 1719 8410
rect 1799 8404 1810 8410
rect 1708 8345 1719 8395
rect 1799 8345 1810 8395
rect 1691 8332 1719 8345
rect 1782 8332 1810 8345
rect 1708 8259 1719 8332
rect 1799 8259 1810 8332
rect 1965 8319 1970 8323
rect 1965 8298 1970 8314
rect 1956 8297 1970 8298
rect 1956 8291 1958 8297
rect 1963 8291 1970 8297
rect 1956 8290 1970 8291
rect 1965 8285 1970 8290
rect 1965 8275 1970 8280
rect 1708 8232 1719 8250
rect 1799 8237 1810 8250
rect 2235 8232 2589 8234
rect 1708 8218 2589 8232
rect 2235 8217 2589 8218
rect 2602 8217 2603 8234
rect 2590 8106 2637 8107
rect 2600 8105 2637 8106
rect 4341 8105 4360 8108
rect 2600 8102 4360 8105
rect 2600 8089 3221 8102
rect 2600 8088 2641 8089
rect 3231 8089 4360 8102
rect 2159 8084 2176 8085
rect 2159 8067 2161 8084
rect 2171 8067 2176 8084
rect 2159 8052 2176 8067
rect 2162 7872 2175 8052
rect 3767 7949 3769 7966
rect 2280 7872 2307 7874
rect 1939 7865 2346 7872
rect 1829 7831 1836 7835
rect 1939 7834 1946 7865
rect 2280 7864 2307 7865
rect 2338 7864 2346 7865
rect 2228 7830 2235 7834
rect 2057 7820 2060 7824
rect 1829 7767 1836 7815
rect 1821 7761 1836 7767
rect 1829 7689 1836 7761
rect 1939 7763 1946 7818
rect 2057 7799 2060 7815
rect 2338 7833 2345 7864
rect 2705 7843 2713 7891
rect 3023 7848 3031 7896
rect 3756 7898 3769 7949
rect 3341 7846 3349 7894
rect 3873 7905 3889 8004
rect 4341 7975 4360 8089
rect 3872 7901 3889 7905
rect 4226 7904 4239 7908
rect 3990 7887 3995 7891
rect 4341 7907 4357 7975
rect 4706 7943 4717 7949
rect 4797 7943 4808 7949
rect 4460 7893 4465 7897
rect 3023 7834 3031 7838
rect 2705 7829 2713 7833
rect 3341 7832 3349 7836
rect 2456 7819 2459 7823
rect 2048 7797 2060 7799
rect 2054 7793 2060 7797
rect 2048 7791 2060 7793
rect 2057 7786 2060 7791
rect 2228 7786 2235 7814
rect 2057 7776 2060 7781
rect 2226 7766 2235 7786
rect 1939 7745 1945 7763
rect 2218 7762 2235 7766
rect 2226 7746 2235 7762
rect 1938 7689 1945 7745
rect 2228 7688 2235 7746
rect 2338 7725 2345 7817
rect 2456 7798 2459 7814
rect 2447 7796 2459 7798
rect 2453 7792 2459 7796
rect 2447 7790 2459 7792
rect 2456 7785 2459 7790
rect 2456 7775 2459 7780
rect 2708 7779 2715 7785
rect 3026 7784 3033 7790
rect 3344 7782 3351 7788
rect 3026 7770 3033 7774
rect 2708 7765 2715 7769
rect 3032 7765 3033 7770
rect 3344 7768 3351 7772
rect 2714 7760 2715 7765
rect 3350 7763 3351 7768
rect 3756 7762 3769 7882
rect 3872 7825 3889 7885
rect 3990 7866 3995 7882
rect 3981 7864 3995 7866
rect 3987 7860 3995 7864
rect 3981 7858 3995 7860
rect 3990 7853 3995 7858
rect 3990 7843 3995 7848
rect 3872 7765 3885 7825
rect 4226 7768 4239 7888
rect 4341 7832 4357 7891
rect 4460 7872 4465 7888
rect 4451 7870 4465 7872
rect 4457 7866 4465 7870
rect 4451 7864 4465 7866
rect 4460 7859 4465 7864
rect 4460 7849 4465 7854
rect 4342 7771 4355 7832
rect 4706 7826 4717 7934
rect 4797 7874 4808 7934
rect 4797 7862 4808 7867
rect 4796 7820 4808 7862
rect 4963 7858 4968 7862
rect 4963 7837 4968 7853
rect 4954 7836 4968 7837
rect 4954 7830 4956 7836
rect 4961 7830 4968 7836
rect 4954 7829 4968 7830
rect 4963 7824 4968 7829
rect 4706 7798 4717 7814
rect 4797 7798 4808 7820
rect 4963 7814 4968 7819
rect 4706 7776 4717 7789
rect 4797 7776 4808 7789
rect 3756 7741 3769 7746
rect 3872 7744 3885 7749
rect 2338 7708 2344 7725
rect 2338 7688 2346 7708
rect 2673 7707 2675 7710
rect 2991 7712 2993 7715
rect 3309 7710 3311 7713
rect 2673 7694 2675 7703
rect 2991 7699 2993 7708
rect 2987 7697 2993 7699
rect 2669 7692 2675 7694
rect 2991 7692 2993 7697
rect 3309 7697 3311 7706
rect 3305 7695 3311 7697
rect 1829 7674 1836 7678
rect 1828 7076 1835 7080
rect 1938 7079 1945 7679
rect 2673 7687 2675 7692
rect 3309 7690 3311 7695
rect 4226 7703 4239 7752
rect 4342 7750 4355 7755
rect 2991 7685 2993 7688
rect 4226 7686 4239 7687
rect 3309 7683 3311 7686
rect 2673 7680 2675 7683
rect 2228 7673 2235 7677
rect 2338 7666 2346 7677
rect 2229 7081 2236 7085
rect 2056 7065 2059 7069
rect 2339 7084 2346 7666
rect 3041 7668 3054 7670
rect 2723 7663 2736 7665
rect 2723 7658 2725 7663
rect 2731 7658 2736 7663
rect 2723 7622 2736 7658
rect 3041 7663 3043 7668
rect 3049 7663 3054 7668
rect 3041 7627 3054 7663
rect 3359 7666 3372 7668
rect 3359 7661 3361 7666
rect 3367 7661 3372 7666
rect 3359 7625 3372 7661
rect 3041 7613 3054 7617
rect 2723 7608 2736 7612
rect 3359 7611 3372 7615
rect 2963 7602 2968 7606
rect 2645 7597 2650 7601
rect 3281 7600 3286 7604
rect 2645 7576 2650 7592
rect 2963 7581 2968 7597
rect 2918 7576 2919 7581
rect 2600 7571 2601 7576
rect 2608 7572 2650 7576
rect 2926 7577 2968 7581
rect 3281 7579 3286 7595
rect 2926 7576 2956 7577
rect 2608 7571 2638 7572
rect 2645 7563 2650 7572
rect 2963 7568 2968 7577
rect 3236 7574 3237 7579
rect 3244 7575 3286 7579
rect 3244 7574 3274 7575
rect 2727 7558 2734 7564
rect 3045 7563 3052 7569
rect 3281 7566 3286 7575
rect 2963 7558 2968 7563
rect 2645 7553 2650 7558
rect 3363 7561 3370 7567
rect 3281 7556 3286 7561
rect 2727 7536 2734 7548
rect 3045 7541 3052 7553
rect 3363 7539 3370 7551
rect 2654 7088 2662 7136
rect 3008 7103 3016 7151
rect 3351 7101 3359 7149
rect 3758 7126 3772 7181
rect 3876 7133 3888 7220
rect 4357 7188 4358 7212
rect 3875 7129 3888 7133
rect 4229 7132 4242 7136
rect 3993 7115 3998 7119
rect 4345 7135 4358 7188
rect 4706 7141 4717 7147
rect 4797 7141 4808 7147
rect 4463 7121 4468 7125
rect 3008 7089 3016 7093
rect 3758 7092 3772 7110
rect 3351 7087 3359 7091
rect 2654 7074 2662 7078
rect 2457 7070 2460 7074
rect 1828 7021 1835 7060
rect 1819 7015 1835 7021
rect 1828 6934 1835 7015
rect 1938 7050 1945 7063
rect 1938 7008 1944 7050
rect 2056 7044 2059 7060
rect 2047 7042 2059 7044
rect 2053 7038 2059 7042
rect 2047 7036 2059 7038
rect 2056 7031 2059 7036
rect 2056 7021 2059 7026
rect 2229 7010 2236 7065
rect 1938 6934 1945 7008
rect 2221 7006 2236 7010
rect 2229 6939 2236 7006
rect 2339 7054 2346 7068
rect 2339 7023 2345 7054
rect 2457 7049 2460 7065
rect 2448 7047 2460 7049
rect 2454 7043 2460 7047
rect 2448 7041 2460 7043
rect 2457 7036 2460 7041
rect 3011 7039 3018 7045
rect 2457 7026 2460 7031
rect 2657 7024 2664 7030
rect 3354 7037 3361 7043
rect 3011 7025 3018 7029
rect 2339 7007 2346 7023
rect 3017 7020 3018 7025
rect 3354 7023 3361 7027
rect 3360 7018 3361 7023
rect 2657 7010 2664 7014
rect 2339 6994 2345 7007
rect 2663 7005 2664 7010
rect 2339 6976 2346 6994
rect 3759 6990 3772 7092
rect 3875 6993 3888 7113
rect 3993 7094 3998 7110
rect 3984 7092 3998 7094
rect 3990 7088 3998 7092
rect 3984 7086 3998 7088
rect 3993 7081 3998 7086
rect 3993 7071 3998 7076
rect 4229 6996 4242 7116
rect 4345 6999 4358 7119
rect 4463 7100 4468 7116
rect 4454 7098 4468 7100
rect 4460 7094 4468 7098
rect 4454 7092 4468 7094
rect 4463 7087 4468 7092
rect 4463 7077 4468 7082
rect 4706 7036 4717 7132
rect 4797 7101 4808 7132
rect 4797 7051 4808 7095
rect 4963 7056 4968 7060
rect 2339 6959 2345 6976
rect 2976 6967 2978 6970
rect 4706 6996 4717 7022
rect 4796 7018 4808 7051
rect 4963 7035 4968 7051
rect 4954 7034 4968 7035
rect 4954 7028 4956 7034
rect 4961 7028 4968 7034
rect 4954 7027 4968 7028
rect 4963 7022 4968 7027
rect 4797 6996 4808 7018
rect 4963 7012 4968 7017
rect 3319 6965 3321 6968
rect 3759 6969 3772 6974
rect 3875 6972 3888 6977
rect 2339 6939 2347 6959
rect 2622 6952 2624 6955
rect 2976 6954 2978 6963
rect 2972 6952 2978 6954
rect 2622 6939 2624 6948
rect 2976 6947 2978 6952
rect 3319 6952 3321 6961
rect 3315 6950 3321 6952
rect 3319 6945 3321 6950
rect 2976 6940 2978 6943
rect 2618 6937 2624 6939
rect 3319 6938 3321 6941
rect 2622 6932 2624 6937
rect 2229 6924 2236 6928
rect 1828 6919 1835 6923
rect 1829 6185 1836 6189
rect 1938 6188 1945 6923
rect 2339 6917 2347 6928
rect 2622 6925 2624 6928
rect 2230 6190 2237 6194
rect 2057 6174 2060 6178
rect 2340 6193 2347 6917
rect 3026 6923 3039 6925
rect 3026 6918 3028 6923
rect 3034 6918 3039 6923
rect 2672 6908 2685 6910
rect 2672 6903 2674 6908
rect 2680 6903 2685 6908
rect 2672 6867 2685 6903
rect 3026 6882 3039 6918
rect 3369 6921 3382 6923
rect 3369 6916 3371 6921
rect 3377 6916 3382 6921
rect 3369 6880 3382 6916
rect 4229 6912 4242 6980
rect 4345 6978 4358 6983
rect 4706 6974 4717 6987
rect 4797 6974 4808 6987
rect 4241 6895 4242 6912
rect 4229 6894 4242 6895
rect 3026 6868 3039 6872
rect 3369 6866 3382 6870
rect 2948 6857 2953 6861
rect 2672 6853 2685 6857
rect 3291 6855 3296 6859
rect 2594 6842 2599 6846
rect 2594 6821 2599 6837
rect 2948 6836 2953 6852
rect 2903 6831 2904 6836
rect 2911 6832 2953 6836
rect 3291 6834 3296 6850
rect 2911 6831 2941 6832
rect 2948 6823 2953 6832
rect 3246 6829 3247 6834
rect 3254 6830 3296 6834
rect 3254 6829 3284 6830
rect 2549 6816 2550 6821
rect 2557 6817 2599 6821
rect 3030 6818 3037 6824
rect 3291 6821 3296 6830
rect 2557 6816 2587 6817
rect 2594 6808 2599 6817
rect 2948 6813 2953 6818
rect 2676 6803 2683 6809
rect 3373 6816 3380 6822
rect 3291 6811 3296 6816
rect 2594 6798 2599 6803
rect 3030 6796 3037 6808
rect 2676 6781 2683 6793
rect 3373 6794 3380 6806
rect 3759 6364 3770 6367
rect 3759 6342 3760 6364
rect 2678 6197 2686 6245
rect 2984 6197 2992 6245
rect 3349 6210 3357 6258
rect 3349 6196 3357 6200
rect 2678 6183 2686 6187
rect 2984 6183 2992 6187
rect 2458 6179 2461 6183
rect 3759 6182 3770 6342
rect 1829 6115 1836 6169
rect 1938 6157 1945 6172
rect 1820 6109 1836 6115
rect 1939 6112 1945 6157
rect 2057 6153 2060 6169
rect 2048 6151 2060 6153
rect 2054 6147 2060 6151
rect 2048 6145 2060 6147
rect 2057 6140 2060 6145
rect 2230 6136 2237 6174
rect 2340 6148 2347 6177
rect 3759 6178 3772 6182
rect 2458 6158 2461 6174
rect 3876 6185 3891 6385
rect 3875 6181 3891 6185
rect 4229 6184 4242 6188
rect 3993 6167 3998 6171
rect 4344 6187 4360 6286
rect 4706 6190 4717 6196
rect 4797 6190 4808 6196
rect 4463 6173 4468 6177
rect 2449 6156 2461 6158
rect 2455 6152 2461 6156
rect 2449 6150 2461 6152
rect 2057 6130 2060 6135
rect 2229 6126 2237 6136
rect 2221 6122 2237 6126
rect 1829 6043 1836 6109
rect 1938 6043 1945 6112
rect 2229 6117 2237 6122
rect 2229 6102 2236 6117
rect 2229 6089 2237 6102
rect 1829 6028 1836 6032
rect 2230 6048 2237 6089
rect 2338 6094 2347 6148
rect 2458 6145 2461 6150
rect 3352 6146 3359 6152
rect 2458 6135 2461 6140
rect 2681 6133 2688 6139
rect 2987 6133 2994 6139
rect 3352 6132 3359 6136
rect 3358 6127 3359 6132
rect 2681 6119 2688 6123
rect 2687 6114 2688 6119
rect 2987 6119 2994 6123
rect 2993 6114 2994 6119
rect 2338 6048 2346 6094
rect 3317 6074 3319 6077
rect 2646 6061 2648 6064
rect 2952 6061 2954 6064
rect 3317 6061 3319 6070
rect 3313 6059 3319 6061
rect 2230 6033 2237 6037
rect 1827 5405 1834 5409
rect 1938 5412 1945 6031
rect 2338 6027 2346 6036
rect 2646 6048 2648 6057
rect 2642 6046 2648 6048
rect 2646 6041 2648 6046
rect 2952 6048 2954 6057
rect 3317 6054 3319 6059
rect 2948 6046 2954 6048
rect 3317 6047 3319 6050
rect 2952 6041 2954 6046
rect 3759 6042 3772 6162
rect 3875 6117 3891 6165
rect 3993 6146 3998 6162
rect 3984 6144 3998 6146
rect 3990 6140 3998 6144
rect 3984 6138 3998 6140
rect 3993 6133 3998 6138
rect 3993 6123 3998 6128
rect 3875 6045 3888 6117
rect 4229 6048 4242 6168
rect 4344 6116 4360 6171
rect 4463 6152 4468 6168
rect 4454 6150 4468 6152
rect 4460 6146 4468 6150
rect 4454 6144 4468 6146
rect 4463 6139 4468 6144
rect 4463 6129 4468 6134
rect 4345 6051 4358 6116
rect 4706 6085 4717 6181
rect 4797 6153 4808 6181
rect 4797 6131 4808 6144
rect 4796 6118 4808 6131
rect 4797 6109 4808 6118
rect 2646 6034 2648 6037
rect 2952 6034 2954 6037
rect 3367 6030 3380 6032
rect 1937 5408 1945 5412
rect 2228 5410 2235 5414
rect 2055 5394 2058 5398
rect 2338 5413 2345 6027
rect 3367 6025 3369 6030
rect 3375 6025 3380 6030
rect 4706 6045 4717 6072
rect 4796 6067 4808 6109
rect 4963 6105 4968 6109
rect 4963 6084 4968 6100
rect 4954 6083 4968 6084
rect 4954 6077 4956 6083
rect 4961 6077 4968 6083
rect 4954 6076 4968 6077
rect 4963 6071 4968 6076
rect 4797 6045 4808 6067
rect 4963 6061 4968 6066
rect 2696 6017 2709 6019
rect 2696 6012 2698 6017
rect 2704 6012 2709 6017
rect 2696 5976 2709 6012
rect 3002 6017 3015 6019
rect 3002 6012 3004 6017
rect 3010 6012 3015 6017
rect 3002 5976 3015 6012
rect 3367 5989 3380 6025
rect 3759 6021 3772 6026
rect 3875 6024 3888 6029
rect 4229 5991 4242 6032
rect 4345 6030 4358 6035
rect 4706 6023 4717 6036
rect 4797 6023 4808 6036
rect 3367 5975 3380 5979
rect 4229 5974 4231 5991
rect 2696 5962 2709 5966
rect 3002 5962 3015 5966
rect 4229 5970 4242 5974
rect 3289 5964 3294 5968
rect 2618 5951 2623 5955
rect 2924 5951 2929 5955
rect 2618 5930 2623 5946
rect 2924 5930 2929 5946
rect 3289 5943 3294 5959
rect 3244 5938 3245 5943
rect 3252 5939 3294 5943
rect 3252 5938 3282 5939
rect 3289 5930 3294 5939
rect 2573 5925 2574 5930
rect 2581 5926 2623 5930
rect 2581 5925 2611 5926
rect 2618 5917 2623 5926
rect 2879 5925 2880 5930
rect 2887 5926 2929 5930
rect 2887 5925 2917 5926
rect 2700 5912 2707 5918
rect 2924 5917 2929 5926
rect 3371 5925 3378 5931
rect 3289 5920 3294 5925
rect 3006 5912 3013 5918
rect 2618 5907 2623 5912
rect 2924 5907 2929 5912
rect 3371 5903 3378 5915
rect 2700 5890 2707 5902
rect 3006 5890 3013 5902
rect 3873 5632 3887 5646
rect 3873 5617 3874 5632
rect 4345 5627 4346 5643
rect 3759 5606 3771 5612
rect 3759 5585 3760 5606
rect 3759 5519 3771 5585
rect 3759 5515 3772 5519
rect 3873 5522 3887 5617
rect 3873 5518 3888 5522
rect 4229 5521 4242 5525
rect 3993 5504 3998 5508
rect 4345 5524 4361 5627
rect 4706 5526 4717 5532
rect 4797 5526 4808 5532
rect 4463 5510 4468 5514
rect 2654 5417 2662 5465
rect 2996 5427 3004 5475
rect 3387 5436 3395 5484
rect 3387 5422 3395 5426
rect 2996 5413 3004 5417
rect 2654 5403 2662 5407
rect 2456 5399 2459 5403
rect 1827 5334 1834 5389
rect 1818 5328 1834 5334
rect 1827 5263 1834 5328
rect 1937 5338 1945 5392
rect 2055 5373 2058 5389
rect 2046 5371 2058 5373
rect 2052 5367 2058 5371
rect 2046 5365 2058 5367
rect 2055 5360 2058 5365
rect 2055 5350 2058 5355
rect 2228 5338 2235 5394
rect 1937 5263 1946 5338
rect 2220 5334 2235 5338
rect 2228 5268 2235 5334
rect 2338 5309 2345 5397
rect 2456 5378 2459 5394
rect 3759 5379 3772 5499
rect 3873 5434 3888 5502
rect 3993 5483 3998 5499
rect 3984 5481 3998 5483
rect 3990 5477 3998 5481
rect 3984 5475 3998 5477
rect 3993 5470 3998 5475
rect 3993 5460 3998 5465
rect 3875 5382 3888 5434
rect 4229 5390 4242 5505
rect 4345 5446 4361 5508
rect 4463 5489 4468 5505
rect 4454 5487 4468 5489
rect 4460 5483 4468 5487
rect 4454 5481 4468 5483
rect 4463 5476 4468 5481
rect 4463 5466 4468 5471
rect 4229 5385 4243 5390
rect 4345 5388 4358 5446
rect 4706 5431 4717 5517
rect 4797 5491 4808 5517
rect 4797 5434 4808 5482
rect 4963 5441 4968 5445
rect 2447 5376 2459 5378
rect 2453 5372 2459 5376
rect 3390 5372 3397 5378
rect 2447 5370 2459 5372
rect 2456 5365 2459 5370
rect 2999 5363 3006 5369
rect 2456 5355 2459 5360
rect 2657 5353 2664 5359
rect 4706 5381 4717 5416
rect 4796 5403 4808 5434
rect 4963 5420 4968 5436
rect 4954 5419 4968 5420
rect 4954 5413 4956 5419
rect 4961 5413 4968 5419
rect 4954 5412 4968 5413
rect 4963 5407 4968 5412
rect 4797 5381 4808 5403
rect 4963 5397 4968 5402
rect 3390 5358 3397 5362
rect 3759 5358 3772 5363
rect 3875 5361 3888 5366
rect 3396 5353 3397 5358
rect 2999 5349 3006 5353
rect 3005 5344 3006 5349
rect 2657 5339 2664 5343
rect 2663 5334 2664 5339
rect 2338 5268 2344 5309
rect 3355 5300 3357 5303
rect 4229 5300 4243 5369
rect 4345 5367 4358 5372
rect 4706 5359 4717 5372
rect 4797 5359 4808 5372
rect 2964 5291 2966 5294
rect 2622 5281 2624 5284
rect 2622 5268 2624 5277
rect 2964 5278 2966 5287
rect 3355 5287 3357 5296
rect 3351 5285 3357 5287
rect 3355 5280 3357 5285
rect 4229 5281 4230 5300
rect 2960 5276 2966 5278
rect 2964 5271 2966 5276
rect 3355 5273 3357 5276
rect 2618 5266 2624 5268
rect 2622 5261 2624 5266
rect 2964 5264 2966 5267
rect 2228 5253 2235 5257
rect 1827 5248 1834 5252
rect 1937 5239 1946 5252
rect 2338 5251 2344 5258
rect 2622 5254 2624 5257
rect 3405 5256 3418 5258
rect 3405 5251 3407 5256
rect 3413 5251 3418 5256
rect 2338 5239 2347 5251
rect 3014 5247 3027 5249
rect 3014 5242 3016 5247
rect 3022 5242 3027 5247
rect 1937 5230 2347 5239
rect 2672 5237 2685 5239
rect 2672 5232 2674 5237
rect 2680 5232 2685 5237
rect 2672 5196 2685 5232
rect 3014 5206 3027 5242
rect 3405 5215 3418 5251
rect 3405 5201 3418 5205
rect 3014 5192 3027 5196
rect 3327 5190 3332 5194
rect 2672 5182 2685 5186
rect 2936 5181 2941 5185
rect 2594 5171 2599 5175
rect 2594 5150 2599 5166
rect 2936 5160 2941 5176
rect 3327 5169 3332 5185
rect 3282 5164 3283 5169
rect 3290 5165 3332 5169
rect 3290 5164 3320 5165
rect 2891 5155 2892 5160
rect 2899 5156 2941 5160
rect 3327 5156 3332 5165
rect 2899 5155 2929 5156
rect 2549 5145 2550 5150
rect 2557 5146 2599 5150
rect 2936 5147 2941 5156
rect 3409 5151 3416 5157
rect 2557 5145 2587 5146
rect 2594 5137 2599 5146
rect 3018 5142 3025 5148
rect 3327 5146 3332 5151
rect 2676 5132 2683 5138
rect 2936 5137 2941 5142
rect 2594 5127 2599 5132
rect 2676 5110 2683 5122
rect 3018 5120 3025 5132
rect 3409 5129 3416 5141
<< polycontact >>
rect 1958 8291 1963 8297
rect 2589 8216 2602 8234
rect 2590 8088 2600 8106
rect 3221 8088 3231 8102
rect 2161 8067 2171 8084
rect 3873 8004 3890 8019
rect 3756 7949 3767 7967
rect 2705 7891 2713 7899
rect 3023 7896 3031 7904
rect 3341 7894 3349 7902
rect 2048 7793 2054 7797
rect 2447 7792 2453 7796
rect 3026 7765 3032 7770
rect 2708 7760 2714 7765
rect 3344 7763 3350 7768
rect 3981 7860 3987 7864
rect 4451 7866 4457 7870
rect 4797 7867 4808 7874
rect 4703 7814 4720 7826
rect 4956 7830 4961 7836
rect 2665 7691 2669 7695
rect 2983 7696 2987 7700
rect 3301 7694 3305 7698
rect 4226 7687 4239 7703
rect 2725 7658 2731 7663
rect 3043 7663 3049 7668
rect 3361 7661 3367 7666
rect 2601 7570 2608 7576
rect 2919 7575 2926 7581
rect 3237 7573 3244 7579
rect 2727 7530 2734 7536
rect 3045 7535 3052 7541
rect 3363 7533 3370 7539
rect 3875 7220 3889 7237
rect 3758 7181 3772 7201
rect 3008 7151 3016 7159
rect 2654 7136 2662 7144
rect 3351 7149 3359 7157
rect 4344 7188 4357 7212
rect 2047 7038 2053 7042
rect 2448 7043 2454 7047
rect 3011 7020 3017 7025
rect 3354 7018 3360 7023
rect 2657 7005 2663 7010
rect 3984 7088 3990 7092
rect 4454 7094 4460 7098
rect 4797 7095 4808 7101
rect 4706 7022 4717 7036
rect 4956 7028 4961 7034
rect 2968 6951 2972 6955
rect 2614 6936 2618 6940
rect 3311 6949 3315 6953
rect 3028 6918 3034 6923
rect 2674 6903 2680 6908
rect 3371 6916 3377 6921
rect 4228 6895 4241 6912
rect 2904 6830 2911 6836
rect 3247 6828 3254 6834
rect 2550 6815 2557 6821
rect 3030 6790 3037 6796
rect 3373 6788 3380 6794
rect 2676 6775 2683 6781
rect 3873 6385 3891 6403
rect 3760 6342 3771 6364
rect 3349 6258 3357 6266
rect 2678 6245 2686 6253
rect 2984 6245 2992 6253
rect 2048 6147 2054 6151
rect 4344 6286 4360 6313
rect 2449 6152 2455 6156
rect 3352 6127 3358 6132
rect 2681 6114 2687 6119
rect 2987 6114 2993 6119
rect 3309 6058 3313 6062
rect 2638 6045 2642 6049
rect 2944 6045 2948 6049
rect 3984 6140 3990 6144
rect 4454 6146 4460 6150
rect 4796 6144 4808 6153
rect 4706 6072 4717 6085
rect 3369 6025 3375 6030
rect 4956 6077 4961 6083
rect 2698 6012 2704 6017
rect 3004 6012 3010 6017
rect 4231 5974 4244 5991
rect 3245 5937 3252 5943
rect 2574 5924 2581 5930
rect 2880 5924 2887 5930
rect 2700 5884 2707 5890
rect 3371 5897 3378 5903
rect 3006 5884 3013 5890
rect 3874 5617 3892 5632
rect 4346 5627 4361 5644
rect 3760 5585 3771 5606
rect 3387 5484 3395 5492
rect 2996 5475 3004 5483
rect 2654 5465 2662 5473
rect 2046 5367 2052 5371
rect 3984 5477 3990 5481
rect 4454 5483 4460 5487
rect 4796 5482 4808 5491
rect 4706 5416 4717 5431
rect 2447 5372 2453 5376
rect 4956 5413 4961 5419
rect 3390 5353 3396 5358
rect 2999 5344 3005 5349
rect 2657 5334 2663 5339
rect 2614 5265 2618 5269
rect 2956 5275 2960 5279
rect 3347 5284 3351 5288
rect 4230 5280 4244 5300
rect 3407 5251 3413 5256
rect 3016 5242 3022 5247
rect 2674 5232 2680 5237
rect 3283 5163 3290 5169
rect 2892 5154 2899 5160
rect 2550 5144 2557 5150
rect 3409 5123 3416 5129
rect 3018 5114 3025 5120
rect 2676 5104 2683 5110
<< metal1 >>
rect 1595 8438 1612 8439
rect 1667 8438 1903 8439
rect 1589 8426 1958 8438
rect 1589 8424 1903 8426
rect 1595 7852 1612 8424
rect 1667 8413 1903 8424
rect 1676 8404 1689 8413
rect 1676 8395 1677 8404
rect 1868 8405 1882 8413
rect 1676 8391 1689 8395
rect 1834 8401 1853 8403
rect 1852 8395 1853 8401
rect 1834 8303 1853 8395
rect 1868 8389 1869 8405
rect 1881 8389 1882 8405
rect 1945 8336 1956 8426
rect 1936 8326 1989 8336
rect 1936 8325 1941 8326
rect 1939 8319 1941 8325
rect 1945 8325 1989 8326
rect 1945 8319 1947 8325
rect 1939 8316 1947 8319
rect 1953 8319 1959 8325
rect 1733 8299 1746 8303
rect 1825 8299 1853 8303
rect 1899 8299 1964 8300
rect 1675 8297 1964 8299
rect 1675 8291 1958 8297
rect 1963 8291 1964 8297
rect 1675 8289 1964 8291
rect 1977 8299 1982 8314
rect 2161 8299 2171 8301
rect 1977 8294 2171 8299
rect 1675 8280 1900 8289
rect 1977 8285 1982 8294
rect 1733 8258 1746 8280
rect 1679 8257 1692 8258
rect 1679 8250 1680 8257
rect 1691 8250 1692 8257
rect 1733 8251 1734 8258
rect 1745 8251 1746 8258
rect 1733 8250 1746 8251
rect 1756 8257 1769 8258
rect 1756 8250 1757 8257
rect 1768 8250 1769 8257
rect 1825 8257 1838 8280
rect 1954 8271 1960 8280
rect 1951 8269 1986 8271
rect 1825 8250 1826 8257
rect 1837 8250 1838 8257
rect 1946 8267 1986 8269
rect 1679 8206 1692 8250
rect 1756 8206 1769 8250
rect 1946 8207 1960 8267
rect 1887 8206 1960 8207
rect 1671 8190 1726 8206
rect 1757 8190 1960 8206
rect 1671 8188 1960 8190
rect 1887 8186 1960 8188
rect 2161 8084 2171 8294
rect 2588 8216 2589 8234
rect 2588 8204 2602 8216
rect 2589 8122 2601 8204
rect 2590 8106 2601 8122
rect 2600 8088 2601 8106
rect 2590 8084 2601 8088
rect 2589 8065 2601 8084
rect 3221 8102 3232 8103
rect 3231 8088 3232 8102
rect 3221 7956 3232 8088
rect 3756 8015 3769 8020
rect 3767 7997 3769 8015
rect 3873 8019 3890 8044
rect 3756 7967 3769 7997
rect 4888 7977 4965 7979
rect 4666 7974 4965 7977
rect 3221 7936 3222 7956
rect 3767 7949 3769 7967
rect 4398 7968 4965 7974
rect 4398 7963 4901 7968
rect 3938 7935 4181 7937
rect 3938 7934 4288 7935
rect 4398 7934 4406 7963
rect 4666 7952 4901 7963
rect 4674 7943 4687 7952
rect 4674 7934 4675 7943
rect 4866 7944 4880 7952
rect 2956 7930 2969 7932
rect 2638 7925 2651 7927
rect 2956 7925 3287 7930
rect 3938 7929 4408 7934
rect 4674 7930 4687 7934
rect 4832 7940 4851 7942
rect 4850 7934 4851 7940
rect 4832 7931 4851 7934
rect 2638 7924 3287 7925
rect 3710 7928 3818 7929
rect 3938 7928 4437 7929
rect 3710 7924 4437 7928
rect 2638 7923 4437 7924
rect 2638 7917 3967 7923
rect 2638 7915 3287 7917
rect 2618 7876 2623 7878
rect 2638 7876 2651 7915
rect 2686 7891 2687 7899
rect 2699 7891 2705 7899
rect 2936 7881 2941 7883
rect 2956 7881 2969 7915
rect 3004 7896 3005 7904
rect 3017 7896 3023 7904
rect 2936 7879 3011 7881
rect 2618 7874 2693 7876
rect 2618 7865 2674 7874
rect 2521 7864 2674 7865
rect 2520 7863 2674 7864
rect 2689 7863 2693 7874
rect 2936 7870 2992 7879
rect 2888 7868 2992 7870
rect 3007 7868 3011 7879
rect 3254 7879 3259 7881
rect 3274 7879 3287 7915
rect 3710 7910 3938 7917
rect 3710 7909 3803 7910
rect 3322 7894 3323 7902
rect 3335 7894 3341 7902
rect 3726 7897 3736 7909
rect 3726 7888 3728 7897
rect 3734 7888 3736 7897
rect 3726 7887 3736 7888
rect 3776 7895 3786 7897
rect 3776 7886 3779 7895
rect 3785 7886 3786 7895
rect 3801 7892 3803 7909
rect 3814 7909 3938 7910
rect 3814 7892 3815 7909
rect 3818 7908 3864 7909
rect 3917 7908 3931 7909
rect 3801 7890 3815 7892
rect 3842 7900 3852 7908
rect 3842 7891 3844 7900
rect 3850 7891 3852 7900
rect 3842 7890 3852 7891
rect 3892 7898 3902 7900
rect 3254 7877 3329 7879
rect 3254 7868 3310 7877
rect 2888 7867 3011 7868
rect 2888 7864 2942 7867
rect 3206 7866 3310 7868
rect 3325 7866 3329 7877
rect 3206 7865 3329 7866
rect 3776 7867 3786 7886
rect 3892 7889 3895 7898
rect 3901 7889 3902 7898
rect 3776 7866 3818 7867
rect 3892 7866 3902 7889
rect 3917 7890 3918 7908
rect 3929 7890 3931 7908
rect 3962 7904 3966 7917
rect 4180 7916 4408 7923
rect 4180 7915 4273 7916
rect 3962 7894 4015 7904
rect 3962 7893 3966 7894
rect 3917 7885 3931 7890
rect 3964 7887 3966 7893
rect 3970 7893 4015 7894
rect 4196 7903 4206 7915
rect 4196 7894 4198 7903
rect 4204 7894 4206 7903
rect 4196 7893 4206 7894
rect 4246 7901 4256 7903
rect 3970 7887 3972 7893
rect 3964 7884 3972 7887
rect 3978 7887 3984 7893
rect 4246 7892 4249 7901
rect 4255 7892 4256 7901
rect 4271 7898 4273 7915
rect 4284 7915 4408 7916
rect 4284 7898 4285 7915
rect 4288 7914 4334 7915
rect 4387 7914 4401 7915
rect 4271 7896 4285 7898
rect 4312 7906 4322 7914
rect 4312 7897 4314 7906
rect 4320 7897 4322 7906
rect 4312 7896 4322 7897
rect 4362 7904 4372 7906
rect 4002 7869 4007 7882
rect 4246 7873 4256 7892
rect 4362 7895 4365 7904
rect 4371 7895 4372 7904
rect 4246 7872 4288 7873
rect 4362 7872 4372 7895
rect 4387 7896 4388 7914
rect 4399 7896 4401 7914
rect 4432 7910 4436 7923
rect 4432 7900 4485 7910
rect 4432 7899 4436 7900
rect 4387 7891 4401 7896
rect 4434 7893 4436 7899
rect 4440 7899 4485 7900
rect 4440 7893 4442 7899
rect 4434 7890 4442 7893
rect 4448 7893 4454 7899
rect 4472 7874 4477 7888
rect 4246 7871 4424 7872
rect 4246 7870 4458 7871
rect 4246 7869 4451 7870
rect 3776 7865 3954 7866
rect 2520 7862 2693 7863
rect 2520 7859 2624 7862
rect 2120 7858 2163 7859
rect 2032 7856 2163 7858
rect 2010 7855 2163 7856
rect 1777 7854 2163 7855
rect 2409 7854 2433 7855
rect 1664 7853 2163 7854
rect 2176 7853 2433 7854
rect 2520 7853 2526 7859
rect 1664 7852 2526 7853
rect 1595 7850 2526 7852
rect 1595 7844 2005 7850
rect 1595 7840 1678 7844
rect 1777 7843 2005 7844
rect 1777 7842 1870 7843
rect 1664 7099 1678 7840
rect 1793 7830 1803 7842
rect 1793 7821 1795 7830
rect 1801 7821 1803 7830
rect 1793 7820 1803 7821
rect 1843 7828 1853 7830
rect 1843 7819 1846 7828
rect 1852 7819 1853 7828
rect 1868 7825 1870 7842
rect 1881 7842 2005 7843
rect 1881 7825 1882 7842
rect 1885 7841 1931 7842
rect 1984 7841 1998 7842
rect 1868 7823 1882 7825
rect 1909 7833 1919 7841
rect 1909 7824 1911 7833
rect 1917 7824 1919 7833
rect 1909 7823 1919 7824
rect 1959 7831 1969 7833
rect 1843 7800 1853 7819
rect 1959 7822 1962 7831
rect 1968 7822 1969 7831
rect 1843 7799 1885 7800
rect 1959 7799 1969 7822
rect 1984 7823 1985 7841
rect 1996 7823 1998 7841
rect 2029 7837 2033 7850
rect 2120 7849 2526 7850
rect 2160 7843 2404 7849
rect 2176 7842 2404 7843
rect 2176 7841 2269 7842
rect 2029 7827 2082 7837
rect 2029 7826 2033 7827
rect 1984 7818 1998 7823
rect 2031 7820 2033 7826
rect 2037 7826 2082 7827
rect 2192 7829 2202 7841
rect 2037 7820 2039 7826
rect 2031 7817 2039 7820
rect 2045 7820 2051 7826
rect 2192 7820 2194 7829
rect 2200 7820 2202 7829
rect 2192 7819 2202 7820
rect 2242 7827 2252 7829
rect 1843 7798 1969 7799
rect 2069 7802 2074 7815
rect 2242 7818 2245 7827
rect 2251 7818 2252 7827
rect 2267 7824 2269 7841
rect 2280 7841 2404 7842
rect 2428 7847 2526 7849
rect 2280 7824 2281 7841
rect 2284 7840 2330 7841
rect 2383 7840 2397 7841
rect 2267 7822 2281 7824
rect 2308 7832 2318 7840
rect 2308 7823 2310 7832
rect 2316 7823 2318 7832
rect 2308 7822 2318 7823
rect 2358 7830 2368 7832
rect 1843 7797 2055 7798
rect 1843 7794 2048 7797
rect 1988 7694 1993 7794
rect 2045 7793 2048 7794
rect 2054 7793 2055 7797
rect 2045 7792 2055 7793
rect 2069 7797 2087 7802
rect 2242 7799 2252 7818
rect 2358 7821 2361 7830
rect 2367 7821 2368 7830
rect 2242 7798 2284 7799
rect 2358 7798 2368 7821
rect 2383 7822 2384 7840
rect 2395 7822 2397 7840
rect 2428 7836 2432 7847
rect 2428 7826 2481 7836
rect 2428 7825 2432 7826
rect 2383 7817 2397 7822
rect 2430 7819 2432 7825
rect 2436 7825 2481 7826
rect 2436 7819 2438 7825
rect 2430 7816 2438 7819
rect 2444 7819 2450 7825
rect 2242 7797 2368 7798
rect 2468 7801 2473 7814
rect 2522 7802 2601 7807
rect 2522 7801 2527 7802
rect 2069 7786 2074 7797
rect 2242 7796 2454 7797
rect 2242 7793 2447 7796
rect 2043 7773 2051 7781
rect 1738 7688 1796 7689
rect 1738 7676 1739 7688
rect 1760 7677 1769 7688
rect 2387 7688 2392 7793
rect 2444 7792 2447 7793
rect 2453 7792 2454 7796
rect 2444 7791 2454 7792
rect 2468 7796 2527 7801
rect 2468 7785 2473 7796
rect 2443 7768 2451 7779
rect 2443 7760 2444 7768
rect 2618 7726 2623 7859
rect 2681 7840 2689 7841
rect 2681 7834 2682 7840
rect 2688 7834 2689 7840
rect 2681 7805 2689 7834
rect 2645 7794 2689 7805
rect 2632 7793 2689 7794
rect 2681 7779 2689 7793
rect 2688 7771 2689 7779
rect 2681 7770 2689 7771
rect 2745 7840 2754 7841
rect 2745 7834 2746 7840
rect 2752 7834 2754 7840
rect 2745 7808 2754 7834
rect 2745 7800 2791 7808
rect 2745 7779 2754 7800
rect 2783 7799 2791 7800
rect 2745 7771 2746 7779
rect 2753 7771 2754 7779
rect 2745 7770 2754 7771
rect 2808 7812 2810 7817
rect 2808 7807 2919 7812
rect 2808 7806 2895 7807
rect 2808 7793 2810 7806
rect 2708 7765 2715 7767
rect 2704 7760 2708 7765
rect 2714 7760 2715 7765
rect 2618 7723 2698 7726
rect 2618 7722 2623 7723
rect 2627 7722 2698 7723
rect 2173 7687 2197 7688
rect 1760 7676 1796 7677
rect 2180 7676 2197 7687
rect 2215 7676 2216 7688
rect 2180 7675 2216 7676
rect 2619 7651 2623 7722
rect 2662 7720 2698 7722
rect 2662 7715 2697 7720
rect 2662 7713 2686 7715
rect 2669 7707 2672 7713
rect 2692 7713 2697 7715
rect 2660 7695 2669 7696
rect 2660 7691 2665 7695
rect 2676 7695 2679 7703
rect 2704 7695 2715 7760
rect 2676 7690 2739 7695
rect 2676 7687 2679 7690
rect 2669 7679 2672 7683
rect 2669 7672 2673 7679
rect 2724 7663 2731 7690
rect 2724 7658 2725 7663
rect 2619 7649 2703 7651
rect 2619 7641 2687 7649
rect 2702 7641 2703 7649
rect 2619 7639 2703 7641
rect 2619 7614 2623 7639
rect 2700 7619 2708 7620
rect 2616 7604 2670 7614
rect 2616 7603 2621 7604
rect 2619 7597 2621 7603
rect 2625 7603 2670 7604
rect 2700 7613 2701 7619
rect 2707 7613 2708 7619
rect 2625 7597 2627 7603
rect 2601 7596 2608 7597
rect 2607 7583 2608 7596
rect 2619 7594 2627 7597
rect 2633 7597 2639 7603
rect 2601 7576 2608 7583
rect 2657 7578 2662 7592
rect 2657 7577 2665 7578
rect 2700 7577 2708 7613
rect 2657 7571 2708 7577
rect 2657 7563 2662 7571
rect 2700 7558 2708 7571
rect 2634 7549 2640 7558
rect 2707 7550 2708 7558
rect 2700 7549 2708 7550
rect 2764 7619 2773 7620
rect 2764 7613 2765 7619
rect 2771 7613 2773 7619
rect 2764 7590 2773 7613
rect 2791 7590 2810 7793
rect 2936 7731 2941 7864
rect 3206 7862 3260 7865
rect 3776 7864 3988 7865
rect 3776 7863 3981 7864
rect 2999 7845 3007 7846
rect 2999 7839 3000 7845
rect 3006 7839 3007 7845
rect 2999 7810 3007 7839
rect 2963 7799 3007 7810
rect 2950 7798 3007 7799
rect 2999 7784 3007 7798
rect 3006 7776 3007 7784
rect 2999 7775 3007 7776
rect 3063 7845 3072 7846
rect 3063 7839 3064 7845
rect 3070 7839 3072 7845
rect 3063 7813 3072 7839
rect 3063 7805 3111 7813
rect 3063 7784 3072 7805
rect 3101 7804 3111 7805
rect 3063 7776 3064 7784
rect 3071 7776 3072 7784
rect 3063 7775 3072 7776
rect 3026 7770 3033 7772
rect 3022 7765 3026 7770
rect 3032 7765 3033 7770
rect 2936 7728 3016 7731
rect 2936 7727 2941 7728
rect 2945 7727 3016 7728
rect 2937 7656 2941 7727
rect 2980 7725 3016 7727
rect 2980 7720 3015 7725
rect 2980 7718 3004 7720
rect 2987 7712 2990 7718
rect 3010 7718 3015 7720
rect 2978 7700 2987 7701
rect 2978 7696 2983 7700
rect 2994 7700 2997 7708
rect 3022 7700 3033 7765
rect 3254 7729 3259 7862
rect 3775 7860 3981 7863
rect 3987 7860 3988 7864
rect 3775 7859 3988 7860
rect 4002 7859 4039 7869
rect 3775 7853 3955 7859
rect 4002 7853 4007 7859
rect 3775 7852 3832 7853
rect 3317 7843 3325 7844
rect 3317 7837 3318 7843
rect 3324 7837 3325 7843
rect 3317 7808 3325 7837
rect 3281 7797 3325 7808
rect 3268 7796 3325 7797
rect 3317 7782 3325 7796
rect 3324 7774 3325 7782
rect 3317 7773 3325 7774
rect 3381 7843 3390 7844
rect 3381 7837 3382 7843
rect 3388 7837 3390 7843
rect 3381 7811 3390 7837
rect 3381 7803 3429 7811
rect 3381 7782 3390 7803
rect 3419 7802 3429 7803
rect 3381 7774 3382 7782
rect 3389 7774 3390 7782
rect 3381 7773 3390 7774
rect 3344 7768 3351 7770
rect 3340 7763 3344 7768
rect 3350 7763 3351 7768
rect 3254 7726 3334 7729
rect 3254 7725 3259 7726
rect 3263 7725 3334 7726
rect 2994 7695 3057 7700
rect 2994 7692 2997 7695
rect 2987 7684 2990 7688
rect 2987 7677 2991 7684
rect 3042 7668 3049 7695
rect 3042 7663 3043 7668
rect 2937 7654 3021 7656
rect 2937 7646 3005 7654
rect 3020 7646 3021 7654
rect 2937 7644 3021 7646
rect 3255 7654 3259 7725
rect 3298 7723 3334 7725
rect 3298 7718 3333 7723
rect 3298 7716 3322 7718
rect 3305 7710 3308 7716
rect 3328 7716 3333 7718
rect 3296 7698 3305 7699
rect 3296 7694 3301 7698
rect 3312 7698 3315 7706
rect 3340 7698 3351 7763
rect 3915 7764 3932 7853
rect 3979 7839 3985 7848
rect 4026 7827 4039 7859
rect 4245 7866 4451 7869
rect 4457 7866 4458 7870
rect 4245 7865 4458 7866
rect 4472 7868 4797 7874
rect 4245 7859 4425 7865
rect 4472 7859 4477 7868
rect 4245 7858 4302 7859
rect 4385 7770 4402 7859
rect 4449 7845 4455 7854
rect 4832 7839 4841 7931
rect 4866 7928 4867 7944
rect 4879 7928 4880 7944
rect 4954 7875 4964 7968
rect 4934 7865 4988 7875
rect 4934 7864 4939 7865
rect 4937 7858 4939 7864
rect 4943 7864 4988 7865
rect 4943 7858 4945 7864
rect 4937 7855 4945 7858
rect 4951 7858 4957 7864
rect 4975 7840 4980 7853
rect 4998 7840 5013 7842
rect 4731 7838 4744 7839
rect 4823 7838 4841 7839
rect 4897 7838 4962 7839
rect 4730 7837 4841 7838
rect 4852 7837 4962 7838
rect 4730 7836 4962 7837
rect 4730 7830 4956 7836
rect 4961 7830 4962 7836
rect 4730 7828 4962 7830
rect 4975 7832 5013 7840
rect 4677 7814 4703 7826
rect 4730 7815 4743 7828
rect 4730 7808 4744 7815
rect 4731 7797 4744 7808
rect 3728 7758 3741 7760
rect 3728 7757 3742 7758
rect 3728 7747 3729 7757
rect 3740 7747 3742 7757
rect 3915 7752 3918 7764
rect 3930 7752 3932 7764
rect 3915 7751 3932 7752
rect 4198 7764 4211 7766
rect 4198 7763 4212 7764
rect 4198 7753 4199 7763
rect 4210 7753 4212 7763
rect 4385 7758 4388 7770
rect 4400 7758 4402 7770
rect 4385 7757 4402 7758
rect 4677 7796 4690 7797
rect 4677 7789 4678 7796
rect 4689 7789 4690 7796
rect 4731 7790 4732 7797
rect 4743 7790 4744 7797
rect 4731 7789 4744 7790
rect 4754 7796 4767 7797
rect 4754 7789 4755 7796
rect 4766 7789 4767 7796
rect 4823 7796 4836 7828
rect 4975 7824 4980 7832
rect 4952 7810 4958 7819
rect 4823 7789 4824 7796
rect 4835 7789 4836 7796
rect 4946 7806 4958 7810
rect 3728 7731 3742 7747
rect 4198 7737 4212 7753
rect 4677 7749 4690 7789
rect 4192 7735 4262 7737
rect 3722 7729 3792 7731
rect 3742 7720 3792 7729
rect 4212 7726 4262 7735
rect 4754 7745 4767 7789
rect 4946 7745 4951 7806
rect 4690 7738 4951 7745
rect 4889 7737 4951 7738
rect 4226 7703 4239 7704
rect 3312 7693 3375 7698
rect 3312 7690 3315 7693
rect 3305 7682 3308 7686
rect 3305 7675 3309 7682
rect 3360 7666 3367 7693
rect 3360 7661 3361 7666
rect 4226 7660 4239 7687
rect 3255 7652 3339 7654
rect 3255 7644 3323 7652
rect 3338 7644 3339 7652
rect 4226 7645 4227 7660
rect 2937 7619 2941 7644
rect 3255 7642 3339 7644
rect 3018 7624 3026 7625
rect 2934 7609 2988 7619
rect 2934 7608 2939 7609
rect 2937 7602 2939 7608
rect 2943 7608 2988 7609
rect 3018 7618 3019 7624
rect 3025 7618 3026 7624
rect 2943 7602 2945 7608
rect 2764 7582 2810 7590
rect 2764 7558 2773 7582
rect 2791 7579 2810 7582
rect 2919 7601 2926 7602
rect 2925 7588 2926 7601
rect 2937 7599 2945 7602
rect 2951 7602 2957 7608
rect 2919 7581 2926 7588
rect 2975 7583 2980 7597
rect 2975 7582 2983 7583
rect 3018 7582 3026 7618
rect 2975 7576 3026 7582
rect 2975 7568 2980 7576
rect 2764 7550 2765 7558
rect 2772 7550 2773 7558
rect 3018 7563 3026 7576
rect 2952 7554 2958 7563
rect 3025 7555 3026 7563
rect 3018 7554 3026 7555
rect 3082 7624 3091 7625
rect 3082 7618 3083 7624
rect 3089 7618 3091 7624
rect 3082 7595 3091 7618
rect 3255 7617 3259 7642
rect 3336 7622 3344 7623
rect 3252 7607 3306 7617
rect 3252 7606 3257 7607
rect 3255 7600 3257 7606
rect 3261 7606 3306 7607
rect 3336 7616 3337 7622
rect 3343 7616 3344 7622
rect 3261 7600 3263 7606
rect 3237 7599 3244 7600
rect 3082 7593 3124 7595
rect 3082 7587 3110 7593
rect 3082 7563 3091 7587
rect 3243 7586 3244 7599
rect 3255 7597 3263 7600
rect 3269 7600 3275 7606
rect 3237 7579 3244 7586
rect 3293 7581 3298 7595
rect 3293 7580 3301 7581
rect 3336 7580 3344 7616
rect 3293 7574 3344 7580
rect 3293 7566 3298 7574
rect 3082 7555 3083 7563
rect 3090 7555 3091 7563
rect 3082 7554 3091 7555
rect 3336 7561 3344 7574
rect 2764 7549 2773 7550
rect 2641 7542 2644 7549
rect 2959 7547 2962 7554
rect 3270 7552 3276 7561
rect 3343 7553 3344 7561
rect 3336 7552 3344 7553
rect 3400 7622 3409 7623
rect 3400 7616 3401 7622
rect 3407 7616 3409 7622
rect 3400 7593 3409 7616
rect 3400 7591 3442 7593
rect 3400 7585 3428 7591
rect 3400 7561 3409 7585
rect 3400 7553 3401 7561
rect 3408 7553 3409 7561
rect 3400 7552 3409 7553
rect 2949 7546 2962 7547
rect 3277 7545 3280 7552
rect 3267 7544 3280 7545
rect 2631 7541 2644 7542
rect 2543 7535 2569 7536
rect 2542 7520 2543 7535
rect 2719 7530 2727 7536
rect 2734 7530 2737 7536
rect 3037 7535 3045 7541
rect 3052 7535 3055 7541
rect 3355 7533 3363 7539
rect 3370 7533 3373 7539
rect 2542 7501 2574 7520
rect 2547 7171 2560 7501
rect 4998 7471 5013 7832
rect 4993 7408 5013 7471
rect 3223 7277 4443 7298
rect 3227 7271 3235 7277
rect 3227 7267 3236 7271
rect 3229 7198 3236 7267
rect 3875 7248 3876 7264
rect 3875 7237 3890 7248
rect 3771 7216 3772 7228
rect 3889 7220 3890 7237
rect 4400 7222 4434 7277
rect 4993 7222 5011 7408
rect 3758 7201 3772 7216
rect 2941 7185 2954 7187
rect 2587 7183 2954 7185
rect 2587 7179 3278 7183
rect 4342 7212 5025 7222
rect 4342 7188 4344 7212
rect 4357 7205 5025 7212
rect 4357 7188 4363 7205
rect 2587 7175 3732 7179
rect 2587 7172 2954 7175
rect 2542 7142 2574 7171
rect 2567 7121 2572 7123
rect 2587 7121 2600 7172
rect 2635 7136 2636 7144
rect 2648 7136 2654 7144
rect 2921 7136 2926 7138
rect 2941 7136 2954 7172
rect 3284 7171 3732 7175
rect 2989 7151 2990 7159
rect 3002 7151 3008 7159
rect 2921 7134 2996 7136
rect 2921 7125 2977 7134
rect 2873 7123 2977 7125
rect 2992 7123 2996 7134
rect 3264 7134 3269 7136
rect 3284 7134 3297 7171
rect 3707 7158 3732 7171
rect 4666 7165 4964 7168
rect 4183 7162 4291 7163
rect 4408 7162 4964 7165
rect 3707 7157 3740 7158
rect 3332 7149 3333 7157
rect 3345 7149 3351 7157
rect 3707 7156 3821 7157
rect 3938 7156 4901 7162
rect 3707 7151 4440 7156
rect 3707 7147 4411 7151
rect 3713 7144 4411 7147
rect 3713 7138 3941 7144
rect 3713 7137 3806 7138
rect 3264 7132 3339 7134
rect 3264 7123 3320 7132
rect 2873 7122 2996 7123
rect 2567 7119 2642 7121
rect 2873 7119 2927 7122
rect 3229 7121 3320 7123
rect 3335 7121 3339 7132
rect 3229 7120 3339 7121
rect 3729 7125 3739 7137
rect 2567 7110 2623 7119
rect 2503 7108 2623 7110
rect 2638 7108 2642 7119
rect 2503 7107 2642 7108
rect 2410 7105 2434 7106
rect 2177 7104 2434 7105
rect 2503 7104 2573 7107
rect 2120 7103 2515 7104
rect 2033 7101 2514 7103
rect 2009 7100 2514 7101
rect 1776 7099 2405 7100
rect 1664 7095 2405 7099
rect 1664 7089 2004 7095
rect 1664 6209 1678 7089
rect 1776 7088 2004 7089
rect 1776 7087 1869 7088
rect 1792 7075 1802 7087
rect 1792 7066 1794 7075
rect 1800 7066 1802 7075
rect 1792 7065 1802 7066
rect 1842 7073 1852 7075
rect 1842 7064 1845 7073
rect 1851 7064 1852 7073
rect 1867 7070 1869 7087
rect 1880 7087 2004 7088
rect 1880 7070 1881 7087
rect 1884 7086 1930 7087
rect 1983 7086 1997 7087
rect 1867 7068 1881 7070
rect 1908 7078 1918 7086
rect 1908 7069 1910 7078
rect 1916 7069 1918 7078
rect 1908 7068 1918 7069
rect 1958 7076 1968 7078
rect 1842 7045 1852 7064
rect 1958 7067 1961 7076
rect 1967 7067 1968 7076
rect 1842 7044 1884 7045
rect 1958 7044 1968 7067
rect 1983 7068 1984 7086
rect 1995 7068 1997 7086
rect 2028 7082 2032 7095
rect 2120 7094 2405 7095
rect 2177 7093 2405 7094
rect 2177 7092 2270 7093
rect 2028 7072 2081 7082
rect 2028 7071 2032 7072
rect 1983 7063 1997 7068
rect 2030 7065 2032 7071
rect 2036 7071 2081 7072
rect 2193 7080 2203 7092
rect 2193 7071 2195 7080
rect 2201 7071 2203 7080
rect 2036 7065 2038 7071
rect 2030 7062 2038 7065
rect 2044 7065 2050 7071
rect 2193 7070 2203 7071
rect 2243 7078 2253 7080
rect 2243 7069 2246 7078
rect 2252 7069 2253 7078
rect 2268 7075 2270 7092
rect 2281 7092 2405 7093
rect 2429 7098 2514 7100
rect 2281 7075 2282 7092
rect 2285 7091 2331 7092
rect 2384 7091 2398 7092
rect 2268 7073 2282 7075
rect 2309 7083 2319 7091
rect 2309 7074 2311 7083
rect 2317 7074 2319 7083
rect 2309 7073 2319 7074
rect 2359 7081 2369 7083
rect 1842 7043 1968 7044
rect 2068 7046 2073 7060
rect 2243 7050 2253 7069
rect 2359 7072 2362 7081
rect 2368 7072 2369 7081
rect 2243 7049 2285 7050
rect 2359 7049 2369 7072
rect 2384 7073 2385 7091
rect 2396 7073 2398 7091
rect 2429 7087 2433 7098
rect 2429 7077 2482 7087
rect 2429 7076 2433 7077
rect 2384 7068 2398 7073
rect 2431 7070 2433 7076
rect 2437 7076 2482 7077
rect 2437 7070 2439 7076
rect 2431 7067 2439 7070
rect 2445 7070 2451 7076
rect 2243 7048 2369 7049
rect 2469 7052 2474 7065
rect 2243 7047 2455 7048
rect 2068 7045 2091 7046
rect 1842 7042 2054 7043
rect 1842 7039 2047 7042
rect 1987 6939 1992 7039
rect 2044 7038 2047 7039
rect 2053 7038 2054 7042
rect 2044 7037 2054 7038
rect 2068 7040 2082 7045
rect 2243 7044 2448 7047
rect 2068 7031 2073 7040
rect 2044 7019 2051 7025
rect 2388 7020 2393 7044
rect 2445 7043 2448 7044
rect 2454 7043 2455 7047
rect 2445 7042 2455 7043
rect 2469 7047 2550 7052
rect 2469 7036 2474 7047
rect 2388 6988 2394 7020
rect 2444 7019 2452 7030
rect 2444 7011 2445 7019
rect 2388 6939 2393 6988
rect 2567 6971 2572 7104
rect 2630 7085 2638 7086
rect 2630 7079 2631 7085
rect 2637 7079 2638 7085
rect 2630 7050 2638 7079
rect 2594 7039 2638 7050
rect 2581 7038 2638 7039
rect 2630 7024 2638 7038
rect 2637 7016 2638 7024
rect 2630 7015 2638 7016
rect 2694 7085 2703 7086
rect 2694 7079 2695 7085
rect 2701 7079 2703 7085
rect 2694 7056 2703 7079
rect 2754 7062 2904 7067
rect 2754 7060 2879 7062
rect 2753 7059 2879 7060
rect 2753 7056 2772 7059
rect 2694 7048 2772 7056
rect 2694 7024 2703 7048
rect 2694 7016 2695 7024
rect 2702 7016 2703 7024
rect 2694 7015 2703 7016
rect 2657 7010 2664 7012
rect 2653 7005 2657 7010
rect 2663 7005 2664 7010
rect 2567 6968 2647 6971
rect 2567 6967 2572 6968
rect 2576 6967 2647 6968
rect 1746 6933 1793 6936
rect 1760 6923 1779 6933
rect 1792 6923 1793 6933
rect 2174 6938 2198 6939
rect 2181 6927 2198 6938
rect 2216 6927 2217 6939
rect 2181 6926 2217 6927
rect 1760 6921 1793 6923
rect 1746 6920 1793 6921
rect 2568 6896 2572 6967
rect 2611 6965 2647 6967
rect 2611 6960 2646 6965
rect 2611 6958 2635 6960
rect 2618 6952 2621 6958
rect 2641 6958 2646 6960
rect 2609 6940 2618 6941
rect 2609 6936 2614 6940
rect 2625 6940 2628 6948
rect 2653 6940 2664 7005
rect 2625 6935 2688 6940
rect 2625 6932 2628 6935
rect 2618 6924 2621 6928
rect 2618 6917 2622 6924
rect 2673 6908 2680 6935
rect 2673 6903 2674 6908
rect 2568 6894 2652 6896
rect 2568 6886 2636 6894
rect 2651 6886 2652 6894
rect 2568 6884 2652 6886
rect 2568 6859 2572 6884
rect 2649 6864 2657 6865
rect 2565 6849 2619 6859
rect 2565 6848 2570 6849
rect 2568 6842 2570 6848
rect 2574 6848 2619 6849
rect 2649 6858 2650 6864
rect 2656 6858 2657 6864
rect 2574 6842 2576 6848
rect 2550 6841 2557 6842
rect 2556 6828 2557 6841
rect 2568 6839 2576 6842
rect 2582 6842 2588 6848
rect 2550 6821 2557 6828
rect 2606 6823 2611 6837
rect 2606 6822 2614 6823
rect 2649 6822 2657 6858
rect 2606 6816 2657 6822
rect 2606 6808 2611 6816
rect 2649 6803 2657 6816
rect 2583 6794 2589 6803
rect 2656 6795 2657 6803
rect 2649 6794 2657 6795
rect 2713 6864 2722 6865
rect 2713 6858 2714 6864
rect 2720 6858 2722 6864
rect 2713 6834 2722 6858
rect 2753 6834 2772 7048
rect 2921 6986 2926 7119
rect 3229 7117 3270 7120
rect 2984 7100 2992 7101
rect 2984 7094 2985 7100
rect 2991 7094 2992 7100
rect 2984 7065 2992 7094
rect 2948 7054 2992 7065
rect 2935 7053 2992 7054
rect 2984 7039 2992 7053
rect 2991 7031 2992 7039
rect 2984 7030 2992 7031
rect 3048 7100 3057 7101
rect 3048 7094 3049 7100
rect 3055 7094 3057 7100
rect 3048 7068 3057 7094
rect 3048 7060 3096 7068
rect 3048 7039 3057 7060
rect 3086 7059 3096 7060
rect 3048 7031 3049 7039
rect 3056 7031 3057 7039
rect 3048 7030 3057 7031
rect 3011 7025 3018 7027
rect 3007 7020 3011 7025
rect 3017 7020 3018 7025
rect 2921 6983 3001 6986
rect 2921 6982 2926 6983
rect 2930 6982 3001 6983
rect 2922 6911 2926 6982
rect 2965 6980 3001 6982
rect 2965 6975 3000 6980
rect 2965 6973 2989 6975
rect 2972 6967 2975 6973
rect 2995 6973 3000 6975
rect 2963 6955 2972 6956
rect 2963 6951 2968 6955
rect 2979 6955 2982 6963
rect 3007 6955 3018 7020
rect 3264 6984 3269 7117
rect 3729 7116 3731 7125
rect 3737 7116 3739 7125
rect 3729 7115 3739 7116
rect 3779 7123 3789 7125
rect 3779 7114 3782 7123
rect 3788 7114 3789 7123
rect 3804 7120 3806 7137
rect 3817 7137 3941 7138
rect 3817 7120 3818 7137
rect 3821 7136 3867 7137
rect 3920 7136 3934 7137
rect 3804 7118 3818 7120
rect 3845 7128 3855 7136
rect 3845 7119 3847 7128
rect 3853 7119 3855 7128
rect 3845 7118 3855 7119
rect 3895 7126 3905 7128
rect 3327 7098 3335 7099
rect 3327 7092 3328 7098
rect 3334 7092 3335 7098
rect 3327 7063 3335 7092
rect 3291 7052 3335 7063
rect 3278 7051 3335 7052
rect 3327 7037 3335 7051
rect 3334 7029 3335 7037
rect 3327 7028 3335 7029
rect 3391 7098 3400 7099
rect 3391 7092 3392 7098
rect 3398 7092 3400 7098
rect 3391 7066 3400 7092
rect 3779 7095 3789 7114
rect 3895 7117 3898 7126
rect 3904 7117 3905 7126
rect 3779 7094 3821 7095
rect 3895 7094 3905 7117
rect 3920 7118 3921 7136
rect 3932 7118 3934 7136
rect 3965 7132 3969 7144
rect 4183 7143 4276 7144
rect 3965 7122 4018 7132
rect 3965 7121 3969 7122
rect 3920 7113 3934 7118
rect 3967 7115 3969 7121
rect 3973 7121 4018 7122
rect 4199 7131 4209 7143
rect 4199 7122 4201 7131
rect 4207 7122 4209 7131
rect 4199 7121 4209 7122
rect 4249 7129 4259 7131
rect 3973 7115 3975 7121
rect 3967 7112 3975 7115
rect 3981 7115 3987 7121
rect 4249 7120 4252 7129
rect 4258 7120 4259 7129
rect 4274 7126 4276 7143
rect 4287 7143 4411 7144
rect 4287 7126 4288 7143
rect 4291 7142 4337 7143
rect 4390 7142 4404 7143
rect 4274 7124 4288 7126
rect 4315 7134 4325 7142
rect 4315 7125 4317 7134
rect 4323 7125 4325 7134
rect 4315 7124 4325 7125
rect 4365 7132 4375 7134
rect 4005 7096 4010 7110
rect 4249 7101 4259 7120
rect 4365 7123 4368 7132
rect 4374 7123 4375 7132
rect 4249 7100 4291 7101
rect 4365 7100 4375 7123
rect 4390 7124 4391 7142
rect 4402 7124 4404 7142
rect 4435 7138 4439 7151
rect 4666 7150 4901 7156
rect 4674 7141 4687 7150
rect 4435 7128 4488 7138
rect 4674 7132 4675 7141
rect 4866 7142 4880 7150
rect 4674 7128 4687 7132
rect 4832 7138 4851 7140
rect 4850 7132 4851 7138
rect 4832 7129 4851 7132
rect 4435 7127 4439 7128
rect 4390 7119 4404 7124
rect 4437 7121 4439 7127
rect 4443 7127 4488 7128
rect 4443 7121 4445 7127
rect 4437 7118 4445 7121
rect 4451 7121 4457 7127
rect 4475 7103 4480 7116
rect 4475 7101 4808 7103
rect 4249 7099 4427 7100
rect 4249 7098 4461 7099
rect 4249 7097 4454 7098
rect 4035 7096 4047 7097
rect 3779 7093 3957 7094
rect 3779 7092 3991 7093
rect 3779 7091 3984 7092
rect 3778 7088 3984 7091
rect 3990 7088 3991 7092
rect 3778 7087 3991 7088
rect 4005 7089 4047 7096
rect 3778 7081 3958 7087
rect 4005 7081 4010 7089
rect 3778 7080 3835 7081
rect 3391 7058 3439 7066
rect 3391 7037 3400 7058
rect 3429 7057 3439 7058
rect 3391 7029 3392 7037
rect 3399 7029 3400 7037
rect 3391 7028 3400 7029
rect 3354 7023 3361 7025
rect 3350 7018 3354 7023
rect 3360 7018 3361 7023
rect 3264 6981 3344 6984
rect 3264 6980 3269 6981
rect 3273 6980 3344 6981
rect 2979 6950 3042 6955
rect 2979 6947 2982 6950
rect 2972 6939 2975 6943
rect 2972 6932 2976 6939
rect 3027 6923 3034 6950
rect 3027 6918 3028 6923
rect 2922 6909 3006 6911
rect 2922 6901 2990 6909
rect 3005 6901 3006 6909
rect 2922 6899 3006 6901
rect 2922 6874 2926 6899
rect 3003 6879 3011 6880
rect 2919 6864 2973 6874
rect 2919 6863 2924 6864
rect 2922 6857 2924 6863
rect 2928 6863 2973 6864
rect 3003 6873 3004 6879
rect 3010 6873 3011 6879
rect 2928 6857 2930 6863
rect 2713 6823 2772 6834
rect 2904 6856 2911 6857
rect 2910 6843 2911 6856
rect 2922 6854 2930 6857
rect 2936 6857 2942 6863
rect 2904 6836 2911 6843
rect 2960 6838 2965 6852
rect 2960 6837 2968 6838
rect 3003 6837 3011 6873
rect 2960 6831 3011 6837
rect 2960 6823 2965 6831
rect 2713 6803 2722 6823
rect 2753 6822 2772 6823
rect 3003 6818 3011 6831
rect 2937 6809 2943 6818
rect 3010 6810 3011 6818
rect 3003 6809 3011 6810
rect 3067 6879 3076 6880
rect 3067 6873 3068 6879
rect 3074 6873 3076 6879
rect 3067 6850 3076 6873
rect 3067 6848 3109 6850
rect 3067 6842 3095 6848
rect 3067 6818 3076 6842
rect 3067 6810 3068 6818
rect 3075 6810 3076 6818
rect 3067 6809 3076 6810
rect 2713 6795 2714 6803
rect 2721 6795 2722 6803
rect 2944 6802 2947 6809
rect 2934 6801 2947 6802
rect 2713 6794 2722 6795
rect 2590 6787 2593 6794
rect 3022 6790 3030 6796
rect 3037 6790 3040 6796
rect 2580 6786 2593 6787
rect 2668 6775 2676 6781
rect 2683 6775 2686 6781
rect 3164 6725 3191 6979
rect 3265 6909 3269 6980
rect 3308 6978 3344 6980
rect 3308 6973 3343 6978
rect 3308 6971 3332 6973
rect 3315 6965 3318 6971
rect 3338 6971 3343 6973
rect 3306 6953 3315 6954
rect 3306 6949 3311 6953
rect 3322 6953 3325 6961
rect 3350 6953 3361 7018
rect 3918 6992 3935 7081
rect 3982 7067 3988 7076
rect 4035 7036 4047 7089
rect 4248 7094 4454 7097
rect 4460 7094 4461 7098
rect 4248 7093 4461 7094
rect 4475 7095 4797 7101
rect 4248 7087 4428 7093
rect 4475 7087 4480 7095
rect 4248 7086 4305 7087
rect 4046 7021 4047 7036
rect 4388 6998 4405 7087
rect 4452 7073 4458 7082
rect 4832 7037 4841 7129
rect 4866 7126 4867 7142
rect 4879 7126 4880 7142
rect 4954 7073 4964 7162
rect 4934 7063 4988 7073
rect 4934 7062 4939 7063
rect 4937 7056 4939 7062
rect 4943 7062 4988 7063
rect 4943 7056 4945 7062
rect 4937 7053 4945 7056
rect 4951 7056 4957 7062
rect 4975 7037 4980 7051
rect 4731 7036 4744 7037
rect 4823 7036 4841 7037
rect 4897 7036 4962 7037
rect 4691 7022 4706 7036
rect 4730 7035 4841 7036
rect 4852 7035 4962 7036
rect 4730 7034 4962 7035
rect 4730 7028 4956 7034
rect 4961 7028 4962 7034
rect 4730 7026 4962 7028
rect 4975 7036 4988 7037
rect 4999 7036 5018 7037
rect 4975 7029 5021 7036
rect 4730 7013 4743 7026
rect 4730 7006 4744 7013
rect 3731 6986 3744 6988
rect 3731 6985 3745 6986
rect 3731 6975 3732 6985
rect 3743 6975 3745 6985
rect 3918 6980 3921 6992
rect 3933 6980 3935 6992
rect 3918 6979 3935 6980
rect 4201 6992 4214 6994
rect 4201 6991 4215 6992
rect 4201 6981 4202 6991
rect 4213 6981 4215 6991
rect 4388 6986 4391 6998
rect 4403 6986 4405 6998
rect 4731 6995 4744 7006
rect 4388 6985 4405 6986
rect 4677 6994 4690 6995
rect 4677 6987 4678 6994
rect 4689 6987 4690 6994
rect 4731 6988 4732 6995
rect 4743 6988 4744 6995
rect 4731 6987 4744 6988
rect 4754 6994 4767 6995
rect 4754 6987 4755 6994
rect 4766 6987 4767 6994
rect 4823 6994 4836 7026
rect 4975 7022 4980 7029
rect 4952 7008 4958 7017
rect 4823 6987 4824 6994
rect 4835 6987 4836 6994
rect 4946 7004 4958 7008
rect 3731 6959 3745 6975
rect 4201 6965 4215 6981
rect 4677 6970 4690 6987
rect 4195 6963 4265 6965
rect 3725 6957 3795 6959
rect 3322 6948 3385 6953
rect 3745 6948 3795 6957
rect 4215 6954 4265 6963
rect 4688 6955 4690 6970
rect 3322 6945 3325 6948
rect 3315 6937 3318 6941
rect 3315 6930 3319 6937
rect 3370 6921 3377 6948
rect 4677 6943 4690 6955
rect 4754 6943 4767 6987
rect 4946 6943 4951 7004
rect 4669 6936 4951 6943
rect 4889 6935 4951 6936
rect 3370 6916 3371 6921
rect 4219 6912 4244 6913
rect 3265 6907 3349 6909
rect 3265 6899 3333 6907
rect 3348 6899 3349 6907
rect 3265 6897 3349 6899
rect 3265 6872 3269 6897
rect 4219 6895 4228 6912
rect 4241 6895 4244 6912
rect 3346 6877 3354 6878
rect 3262 6862 3316 6872
rect 3262 6861 3267 6862
rect 3265 6855 3267 6861
rect 3271 6861 3316 6862
rect 3346 6871 3347 6877
rect 3353 6871 3354 6877
rect 3271 6855 3273 6861
rect 3247 6854 3254 6855
rect 3253 6841 3254 6854
rect 3265 6852 3273 6855
rect 3279 6855 3285 6861
rect 3247 6834 3254 6841
rect 3303 6836 3308 6850
rect 3303 6835 3311 6836
rect 3346 6835 3354 6871
rect 3303 6829 3354 6835
rect 3303 6821 3308 6829
rect 3346 6816 3354 6829
rect 3280 6807 3286 6816
rect 3353 6808 3354 6816
rect 3346 6807 3354 6808
rect 3410 6877 3419 6878
rect 3410 6871 3411 6877
rect 3417 6871 3419 6877
rect 3410 6848 3419 6871
rect 3410 6846 3452 6848
rect 3410 6840 3438 6846
rect 3410 6816 3419 6840
rect 3410 6808 3411 6816
rect 3418 6808 3419 6816
rect 3410 6807 3419 6808
rect 3287 6800 3290 6807
rect 3277 6799 3290 6800
rect 3365 6788 3373 6794
rect 3380 6788 3383 6794
rect 4219 6725 4244 6895
rect 3164 6702 4244 6725
rect 4219 6700 4244 6702
rect 2549 6690 2573 6691
rect 2528 6689 2573 6690
rect 2547 6672 2573 6689
rect 2549 6647 2573 6672
rect 2553 6281 2570 6647
rect 4999 6439 5018 7029
rect 3221 6417 5018 6439
rect 3226 6318 3245 6417
rect 3785 6403 3891 6404
rect 3803 6385 3873 6403
rect 3709 6364 3770 6365
rect 3731 6342 3760 6364
rect 3241 6303 3245 6318
rect 4999 6314 5018 6417
rect 4344 6313 5018 6314
rect 4360 6289 5018 6313
rect 4360 6287 5017 6289
rect 2611 6282 3274 6283
rect 3292 6282 3729 6283
rect 2549 6254 2573 6281
rect 2611 6273 3748 6282
rect 2611 6272 2930 6273
rect 2549 6234 2573 6236
rect 2591 6230 2596 6232
rect 2611 6230 2624 6272
rect 2659 6245 2660 6253
rect 2672 6245 2678 6253
rect 2897 6230 2902 6232
rect 2917 6230 2930 6272
rect 3282 6272 3748 6273
rect 2965 6245 2966 6253
rect 2978 6245 2984 6253
rect 3262 6243 3267 6245
rect 3282 6243 3295 6272
rect 3330 6258 3331 6266
rect 3343 6258 3349 6266
rect 3262 6241 3337 6243
rect 3262 6232 3318 6241
rect 3226 6230 3318 6232
rect 3333 6230 3337 6241
rect 2591 6228 2666 6230
rect 2591 6219 2647 6228
rect 2527 6217 2647 6219
rect 2662 6217 2666 6228
rect 2897 6228 2972 6230
rect 2897 6219 2953 6228
rect 2527 6216 2666 6217
rect 2849 6217 2953 6219
rect 2968 6217 2972 6228
rect 3226 6229 3337 6230
rect 3226 6226 3268 6229
rect 2849 6216 2972 6217
rect 2411 6214 2435 6215
rect 2120 6212 2435 6214
rect 2527 6213 2597 6216
rect 2849 6213 2903 6216
rect 2524 6212 2539 6213
rect 2120 6211 2538 6212
rect 2031 6210 2538 6211
rect 2010 6209 2538 6210
rect 1664 6204 2406 6209
rect 1664 6199 2005 6204
rect 1664 5428 1678 6199
rect 1777 6197 2005 6199
rect 1777 6196 1870 6197
rect 1793 6184 1803 6196
rect 1793 6175 1795 6184
rect 1801 6175 1803 6184
rect 1793 6174 1803 6175
rect 1843 6182 1853 6184
rect 1843 6173 1846 6182
rect 1852 6173 1853 6182
rect 1868 6179 1870 6196
rect 1881 6196 2005 6197
rect 2029 6203 2156 6204
rect 1881 6179 1882 6196
rect 1885 6195 1931 6196
rect 1984 6195 1998 6196
rect 1868 6177 1882 6179
rect 1909 6187 1919 6195
rect 1909 6178 1911 6187
rect 1917 6178 1919 6187
rect 1909 6177 1919 6178
rect 1959 6185 1969 6187
rect 1843 6154 1853 6173
rect 1959 6176 1962 6185
rect 1968 6176 1969 6185
rect 1843 6153 1885 6154
rect 1959 6153 1969 6176
rect 1984 6177 1985 6195
rect 1996 6177 1998 6195
rect 2029 6191 2033 6203
rect 2178 6202 2406 6204
rect 2178 6201 2271 6202
rect 2029 6181 2082 6191
rect 2029 6180 2033 6181
rect 1984 6172 1998 6177
rect 2031 6174 2033 6180
rect 2037 6180 2082 6181
rect 2194 6189 2204 6201
rect 2194 6180 2196 6189
rect 2202 6180 2204 6189
rect 2037 6174 2039 6180
rect 2031 6171 2039 6174
rect 2045 6174 2051 6180
rect 2194 6179 2204 6180
rect 2244 6187 2254 6189
rect 2244 6178 2247 6187
rect 2253 6178 2254 6187
rect 2269 6184 2271 6201
rect 2282 6201 2406 6202
rect 2430 6208 2538 6209
rect 2282 6184 2283 6201
rect 2286 6200 2332 6201
rect 2385 6200 2399 6201
rect 2269 6182 2283 6184
rect 2310 6192 2320 6200
rect 2310 6183 2312 6192
rect 2318 6183 2320 6192
rect 2310 6182 2320 6183
rect 2360 6190 2370 6192
rect 1843 6152 1969 6153
rect 2069 6155 2074 6169
rect 2244 6159 2254 6178
rect 2360 6181 2363 6190
rect 2369 6181 2370 6190
rect 2244 6158 2286 6159
rect 2360 6158 2370 6181
rect 2385 6182 2386 6200
rect 2397 6182 2399 6200
rect 2430 6196 2434 6208
rect 2524 6207 2538 6208
rect 2430 6186 2483 6196
rect 2430 6185 2434 6186
rect 2385 6177 2399 6182
rect 2432 6179 2434 6185
rect 2438 6185 2483 6186
rect 2438 6179 2440 6185
rect 2432 6176 2440 6179
rect 2446 6179 2452 6185
rect 2244 6157 2370 6158
rect 2470 6160 2475 6174
rect 2524 6160 2574 6161
rect 2470 6157 2574 6160
rect 2244 6156 2456 6157
rect 1843 6151 2055 6152
rect 1843 6148 2048 6151
rect 1988 6049 1993 6148
rect 2045 6147 2048 6148
rect 2054 6147 2055 6151
rect 2045 6146 2055 6147
rect 2069 6150 2086 6155
rect 2244 6153 2449 6156
rect 2069 6140 2074 6150
rect 2043 6133 2047 6135
rect 2043 6130 2049 6133
rect 1750 6047 1802 6049
rect 1750 6032 1751 6047
rect 1760 6042 1802 6047
rect 1760 6032 1787 6042
rect 1750 6031 1787 6032
rect 2389 6048 2394 6153
rect 2446 6152 2449 6153
rect 2455 6152 2456 6156
rect 2446 6151 2456 6152
rect 2470 6145 2475 6157
rect 2524 6156 2574 6157
rect 2444 6138 2448 6139
rect 2444 6135 2450 6138
rect 2591 6080 2596 6213
rect 2654 6194 2662 6195
rect 2654 6188 2655 6194
rect 2661 6188 2662 6194
rect 2654 6159 2662 6188
rect 2618 6148 2662 6159
rect 2605 6147 2662 6148
rect 2654 6133 2662 6147
rect 2661 6125 2662 6133
rect 2654 6124 2662 6125
rect 2718 6194 2727 6195
rect 2718 6188 2719 6194
rect 2725 6188 2727 6194
rect 2718 6161 2727 6188
rect 2772 6161 2791 6168
rect 2718 6156 2880 6161
rect 2718 6151 2791 6156
rect 2718 6133 2727 6151
rect 2718 6125 2719 6133
rect 2726 6125 2727 6133
rect 2718 6124 2727 6125
rect 2681 6119 2688 6121
rect 2677 6114 2681 6119
rect 2687 6114 2688 6119
rect 2591 6077 2671 6080
rect 2591 6076 2596 6077
rect 2600 6076 2671 6077
rect 2172 6036 2175 6046
rect 2187 6037 2202 6046
rect 2187 6036 2212 6037
rect 1750 6024 1802 6031
rect 2592 6005 2596 6076
rect 2635 6074 2671 6076
rect 2635 6069 2670 6074
rect 2635 6067 2659 6069
rect 2642 6061 2645 6067
rect 2665 6067 2670 6069
rect 2633 6049 2642 6050
rect 2633 6045 2638 6049
rect 2649 6049 2652 6057
rect 2677 6049 2688 6114
rect 2649 6044 2712 6049
rect 2649 6041 2652 6044
rect 2642 6033 2645 6037
rect 2642 6026 2646 6033
rect 2697 6017 2704 6044
rect 2697 6012 2698 6017
rect 2592 6003 2676 6005
rect 2592 5995 2660 6003
rect 2675 5995 2676 6003
rect 2592 5993 2676 5995
rect 2592 5968 2596 5993
rect 2673 5973 2681 5974
rect 2589 5958 2643 5968
rect 2589 5957 2594 5958
rect 2592 5951 2594 5957
rect 2598 5957 2643 5958
rect 2673 5967 2674 5973
rect 2680 5967 2681 5973
rect 2598 5951 2600 5957
rect 2574 5950 2581 5951
rect 2580 5937 2581 5950
rect 2592 5948 2600 5951
rect 2606 5951 2612 5957
rect 2574 5930 2581 5937
rect 2630 5932 2635 5946
rect 2630 5931 2638 5932
rect 2673 5931 2681 5967
rect 2630 5925 2681 5931
rect 2630 5917 2635 5925
rect 2673 5912 2681 5925
rect 2607 5903 2613 5912
rect 2680 5904 2681 5912
rect 2673 5903 2681 5904
rect 2737 5973 2746 5974
rect 2737 5967 2738 5973
rect 2744 5967 2746 5973
rect 2737 5942 2746 5967
rect 2772 5942 2791 6151
rect 2897 6080 2902 6213
rect 2960 6194 2968 6195
rect 2960 6188 2961 6194
rect 2967 6188 2968 6194
rect 2960 6159 2968 6188
rect 2924 6148 2968 6159
rect 2911 6147 2968 6148
rect 2960 6133 2968 6147
rect 2967 6125 2968 6133
rect 2960 6124 2968 6125
rect 3024 6194 3033 6195
rect 3024 6188 3025 6194
rect 3031 6188 3033 6194
rect 3024 6162 3033 6188
rect 3024 6154 3072 6162
rect 3024 6133 3033 6154
rect 3062 6153 3072 6154
rect 3024 6125 3025 6133
rect 3032 6125 3033 6133
rect 3024 6124 3033 6125
rect 2987 6119 2994 6121
rect 2983 6114 2987 6119
rect 2993 6114 2994 6119
rect 2897 6077 2977 6080
rect 2897 6076 2902 6077
rect 2906 6076 2977 6077
rect 2898 6005 2902 6076
rect 2941 6074 2977 6076
rect 2941 6069 2976 6074
rect 2941 6067 2965 6069
rect 2948 6061 2951 6067
rect 2971 6067 2976 6069
rect 2939 6049 2948 6050
rect 2939 6045 2944 6049
rect 2955 6049 2958 6057
rect 2983 6049 2994 6114
rect 3262 6093 3267 6226
rect 3724 6209 3748 6272
rect 4888 6224 4965 6226
rect 4666 6218 4965 6224
rect 4409 6215 4965 6218
rect 4183 6214 4291 6215
rect 4409 6214 4901 6215
rect 4183 6212 4901 6214
rect 3934 6209 4901 6212
rect 3713 6208 3821 6209
rect 3934 6208 4440 6209
rect 3325 6207 3333 6208
rect 3325 6201 3326 6207
rect 3332 6201 3333 6207
rect 3325 6172 3333 6201
rect 3289 6161 3333 6172
rect 3276 6160 3333 6161
rect 3325 6146 3333 6160
rect 3332 6138 3333 6146
rect 3325 6137 3333 6138
rect 3389 6207 3398 6208
rect 3389 6201 3390 6207
rect 3396 6201 3398 6207
rect 3389 6175 3398 6201
rect 3713 6203 4440 6208
rect 3713 6196 4411 6203
rect 3713 6195 4276 6196
rect 3713 6194 4192 6195
rect 3713 6190 3941 6194
rect 3713 6189 3806 6190
rect 3729 6177 3739 6189
rect 3389 6167 3437 6175
rect 3389 6146 3398 6167
rect 3427 6166 3437 6167
rect 3729 6168 3731 6177
rect 3737 6168 3739 6177
rect 3729 6167 3739 6168
rect 3779 6175 3789 6177
rect 3779 6166 3782 6175
rect 3788 6166 3789 6175
rect 3804 6172 3806 6189
rect 3817 6189 3941 6190
rect 3817 6172 3818 6189
rect 3821 6188 3867 6189
rect 3920 6188 3934 6189
rect 3804 6170 3818 6172
rect 3845 6180 3855 6188
rect 3845 6171 3847 6180
rect 3853 6171 3855 6180
rect 3845 6170 3855 6171
rect 3895 6178 3905 6180
rect 3389 6138 3390 6146
rect 3397 6138 3398 6146
rect 3779 6147 3789 6166
rect 3895 6169 3898 6178
rect 3904 6169 3905 6178
rect 3779 6146 3821 6147
rect 3895 6146 3905 6169
rect 3920 6170 3921 6188
rect 3932 6170 3934 6188
rect 3965 6184 3969 6194
rect 3965 6174 4018 6184
rect 3965 6173 3969 6174
rect 3920 6165 3934 6170
rect 3967 6167 3969 6173
rect 3973 6173 4018 6174
rect 4199 6183 4209 6195
rect 4199 6174 4201 6183
rect 4207 6174 4209 6183
rect 4199 6173 4209 6174
rect 4249 6181 4259 6183
rect 3973 6167 3975 6173
rect 3967 6164 3975 6167
rect 3981 6167 3987 6173
rect 4249 6172 4252 6181
rect 4258 6172 4259 6181
rect 4274 6178 4276 6195
rect 4287 6195 4411 6196
rect 4287 6178 4288 6195
rect 4291 6194 4337 6195
rect 4390 6194 4404 6195
rect 4274 6176 4288 6178
rect 4315 6186 4325 6194
rect 4315 6177 4317 6186
rect 4323 6177 4325 6186
rect 4315 6176 4325 6177
rect 4365 6184 4375 6186
rect 4005 6148 4010 6162
rect 4249 6153 4259 6172
rect 4365 6175 4368 6184
rect 4374 6175 4375 6184
rect 4249 6152 4291 6153
rect 4365 6152 4375 6175
rect 4390 6176 4391 6194
rect 4402 6176 4404 6194
rect 4435 6190 4439 6203
rect 4666 6199 4901 6209
rect 4674 6190 4687 6199
rect 4435 6180 4488 6190
rect 4435 6179 4439 6180
rect 4390 6171 4404 6176
rect 4437 6173 4439 6179
rect 4443 6179 4488 6180
rect 4674 6181 4675 6190
rect 4866 6191 4880 6199
rect 4443 6173 4445 6179
rect 4437 6170 4445 6173
rect 4451 6173 4457 6179
rect 4674 6177 4687 6181
rect 4832 6187 4851 6189
rect 4850 6181 4851 6187
rect 4832 6178 4851 6181
rect 4475 6154 4480 6168
rect 4475 6153 4488 6154
rect 4249 6151 4427 6152
rect 4249 6150 4461 6151
rect 4249 6149 4454 6150
rect 3779 6145 3957 6146
rect 3779 6144 3991 6145
rect 3779 6143 3984 6144
rect 3389 6137 3398 6138
rect 3778 6140 3984 6143
rect 3990 6140 3991 6144
rect 3778 6139 3991 6140
rect 4005 6140 4038 6148
rect 3352 6132 3359 6134
rect 3778 6133 3958 6139
rect 4005 6133 4010 6140
rect 3778 6132 3835 6133
rect 3348 6127 3352 6132
rect 3358 6127 3359 6132
rect 3262 6090 3342 6093
rect 3262 6089 3267 6090
rect 3271 6089 3342 6090
rect 3150 6072 3154 6085
rect 2955 6044 3018 6049
rect 2955 6041 2958 6044
rect 2948 6033 2951 6037
rect 2948 6026 2952 6033
rect 3003 6017 3010 6044
rect 3003 6012 3004 6017
rect 2898 6003 2982 6005
rect 2898 5995 2966 6003
rect 2981 5995 2982 6003
rect 2898 5993 2982 5995
rect 2898 5968 2902 5993
rect 2979 5973 2987 5974
rect 2895 5958 2949 5968
rect 2895 5957 2900 5958
rect 2898 5951 2900 5957
rect 2904 5957 2949 5958
rect 2979 5967 2980 5973
rect 2986 5967 2987 5973
rect 2904 5951 2906 5957
rect 2737 5931 2791 5942
rect 2737 5912 2746 5931
rect 2772 5930 2791 5931
rect 2880 5950 2887 5951
rect 2886 5937 2887 5950
rect 2898 5948 2906 5951
rect 2912 5951 2918 5957
rect 2880 5930 2887 5937
rect 2936 5932 2941 5946
rect 2936 5931 2944 5932
rect 2979 5931 2987 5967
rect 2936 5925 2987 5931
rect 2936 5917 2941 5925
rect 2737 5904 2738 5912
rect 2745 5904 2746 5912
rect 2737 5903 2746 5904
rect 2979 5912 2987 5925
rect 2913 5903 2919 5912
rect 2986 5904 2987 5912
rect 2979 5903 2987 5904
rect 3043 5973 3052 5974
rect 3043 5967 3044 5973
rect 3050 5967 3052 5973
rect 3043 5944 3052 5967
rect 3043 5942 3085 5944
rect 3043 5936 3071 5942
rect 3043 5912 3052 5936
rect 3043 5904 3044 5912
rect 3051 5904 3052 5912
rect 3043 5903 3052 5904
rect 2614 5896 2617 5903
rect 2604 5895 2617 5896
rect 2920 5896 2923 5903
rect 2910 5895 2923 5896
rect 2692 5884 2700 5890
rect 2707 5884 2710 5890
rect 2998 5884 3006 5890
rect 3013 5884 3016 5890
rect 2530 5860 2531 5874
rect 2557 5860 2559 5874
rect 2530 5473 2559 5860
rect 3150 5847 3186 6072
rect 3263 6018 3267 6089
rect 3306 6087 3342 6089
rect 3306 6082 3341 6087
rect 3306 6080 3330 6082
rect 3313 6074 3316 6080
rect 3336 6080 3341 6082
rect 3304 6062 3313 6063
rect 3304 6058 3309 6062
rect 3320 6062 3323 6070
rect 3348 6062 3359 6127
rect 3320 6057 3383 6062
rect 3320 6054 3323 6057
rect 3313 6046 3316 6050
rect 3313 6039 3317 6046
rect 3368 6030 3375 6057
rect 3918 6044 3935 6133
rect 3982 6119 3988 6128
rect 4027 6085 4038 6140
rect 4248 6146 4454 6149
rect 4460 6146 4461 6150
rect 4248 6145 4461 6146
rect 4475 6145 4796 6153
rect 4248 6139 4428 6145
rect 4475 6139 4480 6145
rect 4248 6138 4305 6139
rect 4037 6071 4038 6085
rect 4388 6050 4405 6139
rect 4452 6125 4458 6134
rect 4832 6086 4841 6178
rect 4866 6175 4867 6191
rect 4879 6175 4880 6191
rect 4954 6122 4964 6215
rect 4934 6112 4988 6122
rect 4934 6111 4939 6112
rect 4937 6105 4939 6111
rect 4943 6111 4988 6112
rect 4943 6105 4945 6111
rect 4937 6102 4945 6105
rect 4951 6105 4957 6111
rect 4975 6086 4980 6100
rect 4731 6085 4744 6086
rect 4823 6085 4841 6086
rect 4897 6085 4962 6086
rect 4683 6072 4706 6083
rect 4683 6071 4717 6072
rect 4730 6084 4841 6085
rect 4852 6084 4962 6085
rect 4730 6083 4962 6084
rect 4730 6077 4956 6083
rect 4961 6077 4962 6083
rect 4730 6075 4962 6077
rect 4975 6079 5020 6086
rect 4730 6062 4743 6075
rect 4730 6055 4744 6062
rect 3368 6025 3369 6030
rect 3731 6038 3744 6040
rect 3731 6037 3745 6038
rect 3731 6027 3732 6037
rect 3743 6027 3745 6037
rect 3918 6032 3921 6044
rect 3933 6032 3935 6044
rect 3918 6031 3935 6032
rect 4201 6044 4214 6046
rect 4201 6043 4215 6044
rect 4201 6033 4202 6043
rect 4213 6033 4215 6043
rect 4388 6038 4391 6050
rect 4403 6038 4405 6050
rect 4731 6044 4744 6055
rect 4388 6037 4405 6038
rect 4677 6043 4690 6044
rect 3263 6016 3347 6018
rect 3263 6008 3331 6016
rect 3346 6008 3347 6016
rect 3731 6011 3745 6027
rect 4201 6017 4215 6033
rect 4677 6036 4678 6043
rect 4689 6036 4690 6043
rect 4731 6037 4732 6044
rect 4743 6037 4744 6044
rect 4731 6036 4744 6037
rect 4754 6043 4767 6044
rect 4754 6036 4755 6043
rect 4766 6036 4767 6043
rect 4823 6043 4836 6075
rect 4975 6071 4980 6079
rect 4952 6057 4958 6066
rect 4823 6036 4824 6043
rect 4835 6036 4836 6043
rect 4946 6053 4958 6057
rect 4677 6020 4690 6036
rect 4195 6015 4265 6017
rect 3263 6006 3347 6008
rect 3725 6009 3795 6011
rect 3263 5981 3267 6006
rect 3745 6000 3795 6009
rect 4215 6006 4265 6015
rect 4688 6005 4690 6020
rect 4225 5992 4246 5994
rect 4677 5992 4690 6005
rect 4754 5992 4767 6036
rect 4946 5992 4951 6053
rect 4214 5991 4246 5992
rect 3344 5986 3352 5987
rect 3260 5971 3314 5981
rect 3260 5970 3265 5971
rect 3263 5964 3265 5970
rect 3269 5970 3314 5971
rect 3344 5980 3345 5986
rect 3351 5980 3352 5986
rect 3269 5964 3271 5970
rect 3245 5963 3252 5964
rect 3251 5950 3252 5963
rect 3263 5961 3271 5964
rect 3277 5964 3283 5970
rect 3245 5943 3252 5950
rect 3301 5945 3306 5959
rect 3301 5944 3309 5945
rect 3344 5944 3352 5980
rect 3301 5938 3352 5944
rect 3301 5930 3306 5938
rect 3344 5925 3352 5938
rect 3278 5916 3284 5925
rect 3351 5917 3352 5925
rect 3344 5916 3352 5917
rect 3408 5986 3417 5987
rect 3408 5980 3409 5986
rect 3415 5980 3417 5986
rect 3408 5957 3417 5980
rect 4214 5974 4231 5991
rect 4244 5974 4246 5991
rect 4669 5985 4951 5992
rect 4889 5984 4951 5985
rect 4214 5973 4246 5974
rect 3408 5955 3450 5957
rect 3408 5949 3436 5955
rect 3408 5925 3417 5949
rect 3408 5917 3409 5925
rect 3416 5917 3417 5925
rect 3408 5916 3417 5917
rect 3285 5909 3288 5916
rect 3275 5908 3288 5909
rect 3363 5897 3371 5903
rect 3378 5897 3381 5903
rect 4225 5847 4246 5973
rect 3149 5823 4264 5847
rect 4994 5722 5020 6079
rect 3223 5700 5020 5722
rect 3264 5560 3285 5700
rect 4994 5646 5020 5700
rect 4346 5644 5022 5646
rect 3846 5617 3874 5629
rect 4361 5627 5022 5644
rect 4346 5626 5022 5627
rect 4994 5624 5020 5626
rect 3846 5615 3887 5617
rect 3705 5605 3760 5606
rect 3704 5585 3760 5605
rect 3771 5585 3772 5606
rect 3704 5584 3772 5585
rect 3704 5583 3725 5584
rect 4888 5560 4965 5562
rect 4666 5555 4965 5560
rect 3934 5551 4291 5552
rect 4409 5551 4965 5555
rect 3307 5546 3768 5547
rect 3934 5546 4901 5551
rect 3307 5545 3821 5546
rect 3934 5545 4440 5546
rect 3307 5540 4440 5545
rect 3307 5534 4411 5540
rect 3307 5530 3941 5534
rect 3321 5520 3334 5530
rect 3713 5527 3941 5530
rect 3713 5526 3806 5527
rect 3320 5514 3334 5520
rect 3729 5514 3739 5526
rect 3320 5511 3333 5514
rect 2929 5510 3333 5511
rect 2556 5459 2559 5473
rect 2587 5500 3333 5510
rect 3729 5505 3731 5514
rect 3737 5505 3739 5514
rect 3729 5504 3739 5505
rect 3779 5512 3789 5514
rect 2587 5496 2942 5500
rect 2567 5450 2572 5452
rect 2587 5450 2600 5496
rect 2635 5465 2636 5473
rect 2648 5465 2654 5473
rect 2909 5460 2914 5462
rect 2929 5460 2942 5496
rect 2977 5475 2978 5483
rect 2990 5475 2996 5483
rect 3300 5469 3305 5471
rect 3320 5469 3333 5500
rect 3779 5503 3782 5512
rect 3788 5503 3789 5512
rect 3804 5509 3806 5526
rect 3817 5526 3941 5527
rect 3817 5509 3818 5526
rect 3821 5525 3867 5526
rect 3920 5525 3934 5526
rect 3804 5507 3818 5509
rect 3845 5517 3855 5525
rect 3845 5508 3847 5517
rect 3853 5508 3855 5517
rect 3845 5507 3855 5508
rect 3895 5515 3905 5517
rect 3368 5484 3369 5492
rect 3381 5484 3387 5492
rect 3779 5484 3789 5503
rect 3895 5506 3898 5515
rect 3904 5506 3905 5515
rect 3779 5483 3821 5484
rect 3895 5483 3905 5506
rect 3920 5507 3921 5525
rect 3932 5507 3934 5525
rect 3965 5521 3969 5534
rect 4183 5533 4411 5534
rect 4183 5532 4276 5533
rect 3965 5511 4018 5521
rect 3965 5510 3969 5511
rect 3920 5502 3934 5507
rect 3967 5504 3969 5510
rect 3973 5510 4018 5511
rect 4199 5520 4209 5532
rect 4199 5511 4201 5520
rect 4207 5511 4209 5520
rect 4199 5510 4209 5511
rect 4249 5518 4259 5520
rect 3973 5504 3975 5510
rect 3967 5501 3975 5504
rect 3981 5504 3987 5510
rect 4249 5509 4252 5518
rect 4258 5509 4259 5518
rect 4274 5515 4276 5532
rect 4287 5532 4411 5533
rect 4287 5515 4288 5532
rect 4291 5531 4337 5532
rect 4390 5531 4404 5532
rect 4274 5513 4288 5515
rect 4315 5523 4325 5531
rect 4315 5514 4317 5523
rect 4323 5514 4325 5523
rect 4315 5513 4325 5514
rect 4365 5521 4375 5523
rect 4005 5486 4010 5499
rect 4249 5490 4259 5509
rect 4365 5512 4368 5521
rect 4374 5512 4375 5521
rect 4249 5489 4291 5490
rect 4365 5489 4375 5512
rect 4390 5513 4391 5531
rect 4402 5513 4404 5531
rect 4435 5527 4439 5540
rect 4666 5535 4901 5546
rect 4435 5517 4488 5527
rect 4435 5516 4439 5517
rect 4390 5508 4404 5513
rect 4437 5510 4439 5516
rect 4443 5516 4488 5517
rect 4674 5526 4687 5535
rect 4674 5517 4675 5526
rect 4866 5527 4880 5535
rect 4443 5510 4445 5516
rect 4437 5507 4445 5510
rect 4451 5510 4457 5516
rect 4674 5513 4687 5517
rect 4832 5523 4851 5525
rect 4850 5517 4851 5523
rect 4832 5514 4851 5517
rect 4475 5491 4480 5505
rect 4249 5488 4427 5489
rect 4249 5487 4461 5488
rect 4249 5486 4454 5487
rect 3779 5482 3957 5483
rect 3779 5481 3991 5482
rect 3779 5480 3984 5481
rect 3778 5477 3984 5480
rect 3990 5477 3991 5481
rect 3778 5476 3991 5477
rect 4005 5478 4039 5486
rect 3778 5470 3958 5476
rect 4005 5470 4010 5478
rect 3778 5469 3835 5470
rect 3300 5467 3375 5469
rect 2909 5458 2984 5460
rect 3300 5458 3356 5467
rect 2567 5448 2642 5450
rect 2909 5449 2965 5458
rect 2567 5439 2623 5448
rect 2503 5437 2623 5439
rect 2638 5437 2642 5448
rect 2861 5447 2965 5449
rect 2980 5447 2984 5458
rect 3265 5456 3356 5458
rect 3371 5456 3375 5467
rect 3265 5455 3375 5456
rect 3265 5452 3306 5455
rect 2861 5446 2984 5447
rect 2861 5443 2915 5446
rect 2503 5436 2642 5437
rect 2430 5435 2573 5436
rect 2409 5434 2573 5435
rect 2176 5433 2573 5434
rect 2120 5432 2515 5433
rect 2032 5430 2514 5432
rect 2008 5429 2514 5430
rect 1775 5428 2404 5429
rect 1664 5424 2404 5428
rect 1664 5418 2003 5424
rect 1664 5417 1678 5418
rect 1775 5417 2003 5418
rect 1775 5416 1868 5417
rect 1791 5404 1801 5416
rect 1791 5395 1793 5404
rect 1799 5395 1801 5404
rect 1791 5394 1801 5395
rect 1841 5402 1851 5404
rect 1841 5393 1844 5402
rect 1850 5393 1851 5402
rect 1866 5399 1868 5416
rect 1879 5416 2003 5417
rect 1879 5399 1880 5416
rect 1883 5415 1929 5416
rect 1982 5415 1996 5416
rect 1866 5397 1880 5399
rect 1907 5407 1917 5415
rect 1907 5398 1909 5407
rect 1915 5398 1917 5407
rect 1907 5397 1917 5398
rect 1957 5405 1967 5407
rect 1841 5374 1851 5393
rect 1957 5396 1960 5405
rect 1966 5396 1967 5405
rect 1841 5373 1883 5374
rect 1957 5373 1967 5396
rect 1982 5397 1983 5415
rect 1994 5397 1996 5415
rect 2027 5411 2031 5424
rect 2120 5423 2404 5424
rect 2176 5422 2404 5423
rect 2176 5421 2269 5422
rect 2027 5401 2080 5411
rect 2027 5400 2031 5401
rect 1982 5392 1996 5397
rect 2029 5394 2031 5400
rect 2035 5400 2080 5401
rect 2192 5409 2202 5421
rect 2192 5400 2194 5409
rect 2200 5400 2202 5409
rect 2035 5394 2037 5400
rect 2029 5391 2037 5394
rect 2043 5394 2049 5400
rect 2192 5399 2202 5400
rect 2242 5407 2252 5409
rect 2242 5398 2245 5407
rect 2251 5398 2252 5407
rect 2267 5404 2269 5421
rect 2280 5421 2404 5422
rect 2428 5428 2514 5429
rect 2280 5404 2281 5421
rect 2284 5420 2330 5421
rect 2383 5420 2397 5421
rect 2267 5402 2281 5404
rect 2308 5412 2318 5420
rect 2308 5403 2310 5412
rect 2316 5403 2318 5412
rect 2308 5402 2318 5403
rect 2358 5410 2368 5412
rect 1841 5372 1967 5373
rect 2067 5375 2072 5389
rect 2242 5379 2252 5398
rect 2358 5401 2361 5410
rect 2367 5401 2368 5410
rect 2242 5378 2284 5379
rect 2358 5378 2368 5401
rect 2383 5402 2384 5420
rect 2395 5402 2397 5420
rect 2428 5416 2432 5428
rect 2500 5427 2514 5428
rect 2428 5406 2481 5416
rect 2428 5405 2432 5406
rect 2383 5397 2397 5402
rect 2430 5399 2432 5405
rect 2436 5405 2481 5406
rect 2436 5399 2438 5405
rect 2430 5396 2438 5399
rect 2444 5399 2450 5405
rect 2242 5377 2368 5378
rect 2468 5381 2473 5394
rect 2242 5376 2454 5377
rect 1841 5371 2053 5372
rect 1841 5368 2046 5371
rect 1986 5268 1991 5368
rect 2043 5367 2046 5368
rect 2052 5367 2053 5371
rect 2043 5366 2053 5367
rect 2067 5370 2087 5375
rect 2094 5370 2095 5375
rect 2242 5373 2447 5376
rect 2387 5370 2392 5373
rect 2444 5372 2447 5373
rect 2453 5372 2454 5376
rect 2444 5371 2454 5372
rect 2468 5376 2550 5381
rect 2043 5360 2051 5361
rect 2067 5360 2072 5370
rect 2043 5355 2044 5360
rect 2043 5342 2051 5355
rect 2387 5310 2394 5370
rect 2468 5365 2473 5376
rect 2444 5355 2451 5359
rect 2387 5268 2392 5310
rect 2567 5300 2572 5433
rect 2630 5414 2638 5415
rect 2630 5408 2631 5414
rect 2637 5408 2638 5414
rect 2630 5379 2638 5408
rect 2594 5368 2638 5379
rect 2581 5367 2638 5368
rect 2630 5353 2638 5367
rect 2637 5345 2638 5353
rect 2630 5344 2638 5345
rect 2694 5414 2703 5415
rect 2694 5408 2695 5414
rect 2701 5408 2703 5414
rect 2694 5377 2703 5408
rect 2748 5386 2892 5391
rect 2748 5383 2863 5386
rect 2746 5381 2863 5383
rect 2746 5377 2765 5381
rect 2694 5365 2765 5377
rect 2694 5353 2703 5365
rect 2694 5345 2695 5353
rect 2702 5345 2703 5353
rect 2694 5344 2703 5345
rect 2657 5339 2664 5341
rect 2653 5334 2657 5339
rect 2663 5334 2664 5339
rect 2567 5297 2647 5300
rect 2567 5296 2572 5297
rect 2576 5296 2647 5297
rect 1753 5263 1818 5264
rect 1753 5261 1804 5263
rect 1766 5253 1804 5261
rect 2168 5267 2217 5268
rect 2175 5258 2207 5267
rect 2215 5258 2217 5267
rect 2175 5257 2217 5258
rect 1766 5251 1818 5253
rect 2568 5225 2572 5296
rect 2611 5294 2647 5296
rect 2611 5289 2646 5294
rect 2611 5287 2635 5289
rect 2618 5281 2621 5287
rect 2641 5287 2646 5289
rect 2609 5269 2618 5270
rect 2609 5265 2614 5269
rect 2625 5269 2628 5277
rect 2653 5269 2664 5334
rect 2625 5264 2688 5269
rect 2625 5261 2628 5264
rect 2618 5253 2621 5257
rect 2618 5246 2622 5253
rect 2673 5237 2680 5264
rect 2673 5232 2674 5237
rect 2568 5223 2652 5225
rect 2568 5215 2636 5223
rect 2651 5215 2652 5223
rect 2568 5213 2652 5215
rect 2568 5188 2572 5213
rect 2649 5193 2657 5194
rect 2565 5178 2619 5188
rect 2565 5177 2570 5178
rect 2568 5171 2570 5177
rect 2574 5177 2619 5178
rect 2649 5187 2650 5193
rect 2656 5187 2657 5193
rect 2574 5171 2576 5177
rect 2550 5170 2557 5171
rect 2556 5157 2557 5170
rect 2568 5168 2576 5171
rect 2582 5171 2588 5177
rect 2550 5150 2557 5157
rect 2606 5152 2611 5166
rect 2606 5151 2614 5152
rect 2649 5151 2657 5187
rect 2606 5145 2657 5151
rect 2606 5137 2611 5145
rect 2649 5132 2657 5145
rect 2583 5123 2589 5132
rect 2656 5124 2657 5132
rect 2649 5123 2657 5124
rect 2713 5193 2722 5194
rect 2713 5187 2714 5193
rect 2720 5187 2722 5193
rect 2713 5158 2722 5187
rect 2746 5158 2765 5365
rect 2909 5310 2914 5443
rect 2972 5424 2980 5425
rect 2972 5418 2973 5424
rect 2979 5418 2980 5424
rect 2972 5389 2980 5418
rect 2936 5378 2980 5389
rect 2923 5377 2980 5378
rect 2972 5363 2980 5377
rect 2979 5355 2980 5363
rect 2972 5354 2980 5355
rect 3036 5424 3045 5425
rect 3036 5418 3037 5424
rect 3043 5418 3045 5424
rect 3036 5392 3045 5418
rect 3036 5384 3084 5392
rect 3036 5363 3045 5384
rect 3074 5383 3084 5384
rect 3036 5355 3037 5363
rect 3044 5355 3045 5363
rect 3036 5354 3045 5355
rect 2999 5349 3006 5351
rect 2995 5344 2999 5349
rect 3005 5344 3006 5349
rect 2909 5307 2989 5310
rect 2909 5306 2914 5307
rect 2918 5306 2989 5307
rect 2910 5235 2914 5306
rect 2953 5304 2989 5306
rect 2953 5299 2988 5304
rect 2953 5297 2977 5299
rect 2960 5291 2963 5297
rect 2983 5297 2988 5299
rect 2951 5279 2960 5280
rect 2951 5275 2956 5279
rect 2967 5279 2970 5287
rect 2995 5279 3006 5344
rect 3300 5319 3305 5452
rect 3363 5433 3371 5434
rect 3363 5427 3364 5433
rect 3370 5427 3371 5433
rect 3363 5398 3371 5427
rect 3327 5387 3371 5398
rect 3314 5386 3371 5387
rect 3363 5372 3371 5386
rect 3370 5364 3371 5372
rect 3363 5363 3371 5364
rect 3427 5433 3436 5434
rect 3427 5427 3428 5433
rect 3434 5427 3436 5433
rect 3427 5401 3436 5427
rect 3427 5393 3475 5401
rect 3427 5372 3436 5393
rect 3465 5392 3475 5393
rect 3918 5381 3935 5470
rect 3982 5456 3988 5465
rect 4031 5429 4039 5478
rect 4248 5483 4454 5486
rect 4460 5483 4461 5487
rect 4248 5482 4461 5483
rect 4475 5483 4796 5491
rect 4248 5476 4428 5482
rect 4475 5476 4480 5483
rect 4248 5475 4305 5476
rect 4037 5416 4039 5429
rect 4388 5387 4405 5476
rect 4452 5462 4458 5471
rect 4668 5428 4706 5429
rect 4686 5416 4706 5428
rect 4832 5422 4841 5514
rect 4866 5511 4867 5527
rect 4879 5511 4880 5527
rect 4954 5458 4964 5551
rect 4934 5448 4988 5458
rect 4934 5447 4939 5448
rect 4937 5441 4939 5447
rect 4943 5447 4988 5448
rect 4943 5441 4945 5447
rect 4937 5438 4945 5441
rect 4951 5441 4957 5447
rect 4975 5422 4980 5436
rect 4731 5421 4744 5422
rect 4823 5421 4841 5422
rect 4897 5421 4962 5422
rect 4686 5414 4717 5416
rect 4730 5420 4841 5421
rect 4852 5420 4962 5421
rect 4730 5419 4962 5420
rect 4730 5413 4956 5419
rect 4961 5413 4962 5419
rect 4730 5411 4962 5413
rect 4975 5419 4988 5422
rect 4730 5398 4743 5411
rect 4730 5391 4744 5398
rect 3427 5364 3428 5372
rect 3435 5364 3436 5372
rect 3427 5363 3436 5364
rect 3731 5375 3744 5377
rect 3731 5374 3745 5375
rect 3731 5364 3732 5374
rect 3743 5364 3745 5374
rect 3918 5369 3921 5381
rect 3933 5369 3935 5381
rect 3918 5368 3935 5369
rect 4201 5381 4214 5383
rect 4201 5380 4215 5381
rect 4201 5370 4202 5380
rect 4213 5370 4215 5380
rect 4388 5375 4391 5387
rect 4403 5375 4405 5387
rect 4731 5380 4744 5391
rect 4388 5374 4405 5375
rect 4677 5379 4690 5380
rect 3390 5358 3397 5360
rect 3386 5353 3390 5358
rect 3396 5353 3397 5358
rect 3300 5316 3380 5319
rect 3300 5315 3305 5316
rect 3309 5315 3380 5316
rect 3185 5299 3186 5312
rect 2967 5274 3030 5279
rect 2967 5271 2970 5274
rect 2960 5263 2963 5267
rect 2960 5256 2964 5263
rect 3015 5247 3022 5274
rect 3015 5242 3016 5247
rect 2910 5233 2994 5235
rect 2910 5225 2978 5233
rect 2993 5225 2994 5233
rect 2910 5223 2994 5225
rect 2910 5198 2914 5223
rect 2991 5203 2999 5204
rect 2907 5188 2961 5198
rect 2907 5187 2912 5188
rect 2910 5181 2912 5187
rect 2916 5187 2961 5188
rect 2991 5197 2992 5203
rect 2998 5197 2999 5203
rect 2916 5181 2918 5187
rect 2713 5146 2765 5158
rect 2892 5180 2899 5181
rect 2898 5167 2899 5180
rect 2910 5178 2918 5181
rect 2924 5181 2930 5187
rect 2892 5160 2899 5167
rect 2948 5162 2953 5176
rect 2948 5161 2956 5162
rect 2991 5161 2999 5197
rect 2948 5155 2999 5161
rect 2948 5147 2953 5155
rect 2713 5132 2722 5146
rect 2746 5145 2765 5146
rect 2991 5142 2999 5155
rect 2925 5133 2931 5142
rect 2998 5134 2999 5142
rect 2991 5133 2999 5134
rect 3055 5203 3064 5204
rect 3055 5197 3056 5203
rect 3062 5197 3064 5203
rect 3055 5174 3064 5197
rect 3055 5172 3097 5174
rect 3055 5166 3083 5172
rect 3055 5142 3064 5166
rect 3055 5134 3056 5142
rect 3063 5134 3064 5142
rect 3055 5133 3064 5134
rect 2713 5124 2714 5132
rect 2721 5124 2722 5132
rect 2932 5126 2935 5133
rect 2922 5125 2935 5126
rect 2713 5123 2722 5124
rect 2590 5116 2593 5123
rect 2580 5115 2593 5116
rect 3010 5114 3018 5120
rect 3025 5114 3028 5120
rect 2668 5104 2676 5110
rect 2683 5104 2686 5110
rect 3185 5015 3221 5299
rect 3301 5244 3305 5315
rect 3344 5313 3380 5315
rect 3344 5308 3379 5313
rect 3344 5306 3368 5308
rect 3351 5300 3354 5306
rect 3374 5306 3379 5308
rect 3342 5288 3351 5289
rect 3342 5284 3347 5288
rect 3358 5288 3361 5296
rect 3386 5288 3397 5353
rect 3731 5348 3745 5364
rect 4201 5354 4215 5370
rect 4677 5372 4678 5379
rect 4689 5372 4690 5379
rect 4731 5373 4732 5380
rect 4743 5373 4744 5380
rect 4731 5372 4744 5373
rect 4754 5379 4767 5380
rect 4754 5372 4755 5379
rect 4766 5372 4767 5379
rect 4823 5379 4836 5411
rect 4975 5407 4980 5419
rect 4952 5393 4958 5402
rect 4823 5372 4824 5379
rect 4835 5372 4836 5379
rect 4946 5389 4958 5393
rect 4677 5358 4690 5372
rect 4195 5352 4265 5354
rect 3725 5346 3795 5348
rect 3745 5337 3795 5346
rect 4215 5343 4265 5352
rect 4688 5343 4690 5358
rect 4677 5328 4690 5343
rect 4754 5328 4767 5372
rect 4946 5328 4951 5389
rect 4669 5320 4951 5328
rect 3358 5283 3421 5288
rect 3358 5280 3361 5283
rect 3351 5272 3354 5276
rect 3351 5265 3355 5272
rect 3406 5256 3413 5283
rect 4229 5280 4230 5300
rect 4229 5275 4244 5280
rect 4215 5274 4248 5275
rect 3406 5251 3407 5256
rect 4211 5256 4248 5274
rect 3301 5242 3385 5244
rect 3301 5234 3369 5242
rect 3384 5234 3385 5242
rect 3301 5232 3385 5234
rect 3301 5207 3305 5232
rect 3382 5212 3390 5213
rect 3298 5197 3352 5207
rect 3298 5196 3303 5197
rect 3301 5190 3303 5196
rect 3307 5196 3352 5197
rect 3382 5206 3383 5212
rect 3389 5206 3390 5212
rect 3307 5190 3309 5196
rect 3283 5189 3290 5190
rect 3289 5176 3290 5189
rect 3301 5187 3309 5190
rect 3315 5190 3321 5196
rect 3283 5169 3290 5176
rect 3339 5171 3344 5185
rect 3339 5170 3347 5171
rect 3382 5170 3390 5206
rect 3339 5164 3390 5170
rect 3339 5156 3344 5164
rect 3382 5151 3390 5164
rect 3316 5142 3322 5151
rect 3389 5143 3390 5151
rect 3382 5142 3390 5143
rect 3446 5212 3455 5213
rect 3446 5206 3447 5212
rect 3453 5206 3455 5212
rect 3446 5183 3455 5206
rect 3446 5181 3488 5183
rect 3446 5175 3474 5181
rect 3446 5151 3455 5175
rect 3446 5143 3447 5151
rect 3454 5143 3455 5151
rect 3446 5142 3455 5143
rect 3323 5135 3326 5142
rect 3313 5134 3326 5135
rect 3401 5123 3409 5129
rect 3416 5123 3419 5129
rect 4211 5015 4247 5256
rect 3185 4998 4247 5015
rect 3185 4995 4237 4998
<< m2contact >>
rect 1726 8190 1757 8206
rect 2589 8041 2602 8065
rect 3873 8044 3889 8069
rect 2601 7802 2610 7807
rect 2043 7764 2051 7773
rect 1739 7676 1760 7688
rect 2444 7760 2451 7768
rect 2632 7794 2645 7805
rect 2791 7793 2808 7817
rect 2919 7807 2928 7812
rect 2173 7675 2180 7687
rect 2662 7671 2669 7679
rect 2601 7583 2607 7596
rect 2950 7799 2963 7810
rect 3111 7804 3123 7813
rect 3268 7797 3281 7808
rect 3429 7802 3441 7811
rect 2980 7676 2987 7684
rect 3975 7830 3986 7839
rect 4445 7836 4456 7845
rect 3298 7674 3305 7682
rect 2919 7588 2925 7601
rect 3110 7586 3124 7593
rect 3237 7586 3243 7599
rect 2631 7542 2641 7549
rect 2949 7547 2959 7554
rect 3428 7584 3442 7591
rect 3267 7545 3277 7552
rect 3876 7248 3890 7265
rect 2044 7013 2051 7019
rect 2550 7047 2559 7052
rect 2445 7011 2452 7019
rect 2581 7039 2594 7050
rect 2904 7062 2913 7067
rect 1746 6921 1760 6933
rect 2174 6926 2181 6938
rect 2611 6916 2618 6924
rect 2550 6828 2556 6841
rect 2935 7054 2948 7065
rect 3096 7059 3108 7068
rect 3278 7052 3291 7063
rect 3439 7057 3451 7066
rect 2965 6931 2972 6939
rect 2904 6843 2910 6856
rect 3095 6841 3109 6848
rect 2934 6802 2944 6809
rect 2580 6787 2590 6794
rect 3978 7058 3989 7067
rect 4448 7064 4459 7073
rect 3308 6929 3315 6937
rect 3247 6841 3253 6854
rect 3438 6839 3452 6846
rect 3277 6800 3287 6807
rect 3785 6385 3803 6403
rect 2043 6123 2049 6130
rect 1751 6032 1760 6047
rect 2574 6156 2583 6161
rect 2444 6129 2451 6135
rect 2605 6148 2618 6159
rect 2880 6156 2889 6161
rect 2175 6036 2187 6046
rect 2635 6025 2642 6033
rect 2574 5937 2580 5950
rect 2911 6148 2924 6159
rect 3072 6153 3084 6162
rect 3276 6161 3289 6172
rect 3437 6166 3449 6175
rect 2941 6025 2948 6033
rect 2880 5937 2886 5950
rect 3071 5935 3085 5942
rect 2604 5896 2614 5903
rect 2910 5896 2920 5903
rect 3306 6038 3313 6046
rect 3978 6110 3989 6119
rect 4448 6116 4459 6125
rect 3245 5950 3251 5963
rect 3436 5948 3450 5955
rect 3275 5909 3285 5916
rect 3828 5615 3846 5630
rect 2550 5376 2559 5381
rect 2043 5329 2051 5342
rect 2444 5338 2451 5355
rect 2581 5368 2594 5379
rect 2892 5386 2901 5391
rect 1752 5251 1766 5261
rect 2167 5256 2175 5267
rect 2611 5245 2618 5253
rect 2550 5157 2556 5170
rect 2923 5378 2936 5389
rect 3084 5383 3096 5392
rect 3314 5387 3327 5398
rect 3475 5392 3487 5401
rect 3978 5447 3989 5456
rect 4448 5453 4459 5462
rect 2953 5255 2960 5263
rect 2892 5167 2898 5180
rect 3083 5165 3097 5172
rect 2922 5126 2932 5133
rect 2580 5116 2590 5123
rect 3344 5264 3351 5272
rect 3283 5176 3289 5189
rect 3474 5174 3488 5181
rect 3313 5135 3323 5142
<< metal2 >>
rect 1724 8206 1755 8207
rect 1724 8190 1726 8206
rect 1724 7725 1755 8190
rect 2588 8041 2589 8065
rect 2786 8045 3873 8068
rect 2602 8041 2603 8042
rect 2588 8023 2603 8041
rect 2589 7900 2603 8023
rect 2788 8022 2815 8045
rect 2589 7888 2603 7890
rect 2788 7886 2812 8022
rect 2791 7817 2811 7886
rect 2610 7802 2632 7805
rect 2601 7794 2632 7802
rect 2645 7794 2646 7805
rect 2043 7726 2051 7764
rect 2444 7734 2451 7760
rect 2172 7733 2451 7734
rect 2160 7729 2451 7733
rect 2158 7726 2179 7729
rect 2043 7725 2179 7726
rect 1723 7719 2179 7725
rect 1723 7718 2052 7719
rect 1723 7716 1787 7718
rect 1723 7690 1733 7716
rect 2172 7710 2179 7719
rect 2172 7690 2180 7710
rect 1601 7688 1760 7690
rect 1601 7677 1739 7688
rect 1601 6934 1608 7677
rect 2173 7687 2180 7690
rect 2442 7654 2451 7729
rect 2444 7547 2451 7654
rect 2601 7596 2608 7794
rect 2808 7793 2811 7817
rect 3974 7830 3975 7839
rect 3111 7813 3124 7816
rect 2928 7807 2950 7810
rect 2919 7799 2950 7807
rect 2963 7799 2964 7810
rect 3123 7804 3124 7813
rect 3429 7811 3442 7814
rect 2627 7671 2662 7679
rect 2627 7614 2631 7671
rect 2607 7583 2608 7596
rect 2624 7549 2631 7614
rect 2919 7601 2926 7799
rect 3111 7749 3124 7804
rect 3237 7797 3268 7808
rect 3281 7797 3282 7808
rect 3441 7802 3442 7811
rect 3237 7749 3244 7797
rect 3111 7743 3244 7749
rect 2945 7676 2980 7684
rect 2945 7619 2949 7676
rect 2925 7588 2926 7601
rect 2942 7554 2949 7619
rect 3111 7593 3124 7743
rect 3237 7659 3244 7743
rect 3237 7599 3244 7645
rect 3263 7674 3298 7682
rect 3263 7617 3267 7674
rect 3243 7586 3244 7599
rect 2921 7552 2935 7553
rect 2940 7552 2949 7554
rect 2601 7547 2615 7548
rect 2622 7547 2631 7549
rect 2444 7542 2631 7547
rect 2888 7547 2949 7552
rect 3260 7552 3267 7617
rect 3429 7591 3442 7802
rect 3974 7735 3986 7830
rect 4444 7836 4445 7845
rect 4444 7749 4456 7836
rect 4444 7738 4669 7749
rect 4262 7737 4669 7738
rect 4139 7735 4214 7736
rect 3974 7732 4192 7735
rect 3792 7731 4192 7732
rect 3669 7729 3744 7730
rect 3669 7720 3722 7729
rect 3742 7720 3744 7729
rect 3812 7726 4192 7731
rect 4212 7726 4214 7735
rect 4282 7736 4669 7737
rect 4282 7726 4456 7736
rect 3812 7720 4140 7726
rect 3235 7550 3249 7551
rect 3258 7550 3267 7552
rect 2888 7546 2959 7547
rect 2444 7541 2641 7542
rect 2601 7518 2615 7541
rect 2921 7518 2935 7546
rect 3218 7545 3267 7550
rect 3218 7544 3277 7545
rect 3235 7518 3249 7544
rect 3672 7518 3682 7720
rect 2599 7508 3685 7518
rect 3255 7504 3685 7508
rect 2904 7248 3876 7263
rect 3890 7248 3891 7263
rect 2904 7067 2910 7248
rect 3096 7068 3109 7071
rect 2913 7062 2935 7065
rect 2904 7054 2935 7062
rect 2948 7054 2949 7065
rect 3108 7059 3109 7068
rect 3439 7066 3452 7069
rect 2559 7047 2581 7050
rect 2550 7039 2581 7047
rect 2594 7039 2595 7050
rect 2044 6984 2051 7013
rect 2445 7010 2452 7011
rect 2444 6985 2452 7010
rect 2173 6984 2452 6985
rect 1734 6980 1783 6981
rect 2044 6980 2452 6984
rect 1734 6977 2180 6980
rect 1734 6975 2051 6977
rect 1734 6972 1783 6975
rect 1734 6934 1745 6972
rect 2173 6961 2180 6977
rect 2173 6941 2181 6961
rect 2174 6938 2181 6941
rect 1601 6933 1761 6934
rect 1601 6921 1746 6933
rect 1760 6921 1761 6933
rect 1601 6046 1608 6921
rect 2443 6794 2452 6980
rect 2550 6841 2557 7039
rect 2576 6916 2611 6924
rect 2576 6859 2580 6916
rect 2556 6828 2557 6841
rect 2573 6794 2580 6859
rect 2904 6856 2911 7054
rect 3096 6991 3109 7059
rect 3256 7058 3278 7063
rect 3247 7052 3278 7058
rect 3291 7052 3292 7063
rect 3451 7057 3452 7066
rect 3096 6979 3162 6991
rect 3247 6991 3254 7052
rect 3191 6979 3254 6991
rect 2930 6931 2965 6939
rect 2930 6874 2934 6931
rect 2910 6843 2911 6856
rect 2927 6809 2934 6874
rect 3096 6848 3109 6979
rect 3247 6854 3254 6979
rect 3273 6929 3308 6937
rect 3273 6872 3277 6929
rect 3253 6841 3254 6854
rect 2925 6807 2934 6809
rect 2873 6802 2934 6807
rect 3270 6807 3277 6872
rect 3439 6911 3452 7057
rect 3977 7058 3978 7067
rect 3977 6963 3989 7058
rect 4447 7064 4448 7073
rect 4447 6970 4459 7064
rect 4447 6966 4677 6970
rect 4265 6965 4677 6966
rect 4142 6963 4217 6964
rect 3451 6895 3452 6911
rect 3439 6846 3452 6895
rect 3669 6958 3681 6962
rect 3977 6960 4195 6963
rect 3795 6959 4195 6960
rect 3669 6957 3747 6958
rect 3669 6948 3725 6957
rect 3745 6948 3747 6957
rect 3815 6955 4195 6959
rect 3815 6948 3989 6955
rect 4142 6954 4195 6955
rect 4215 6954 4217 6963
rect 4285 6957 4677 6965
rect 4285 6954 4459 6957
rect 4688 6957 4691 6970
rect 3669 6861 3681 6948
rect 3268 6805 3277 6807
rect 2873 6801 2944 6802
rect 2443 6792 2515 6794
rect 2571 6792 2580 6794
rect 2443 6787 2580 6792
rect 2443 6786 2452 6787
rect 2503 6786 2590 6787
rect 2562 6755 2573 6786
rect 2899 6755 2913 6801
rect 3229 6800 3277 6805
rect 3229 6799 3287 6800
rect 3243 6760 3262 6799
rect 3670 6760 3680 6861
rect 3243 6755 3682 6760
rect 2562 6740 3682 6755
rect 2565 6739 3682 6740
rect 3259 6738 3682 6739
rect 2879 6402 3785 6403
rect 2878 6386 3785 6402
rect 2878 6161 2889 6386
rect 3437 6175 3450 6178
rect 3255 6167 3276 6172
rect 2583 6156 2605 6159
rect 2574 6148 2605 6156
rect 2618 6148 2619 6159
rect 2878 6156 2880 6161
rect 3072 6162 3085 6165
rect 2889 6156 2911 6159
rect 2878 6148 2911 6156
rect 2924 6148 2925 6159
rect 3084 6153 3085 6162
rect 2043 6101 2049 6123
rect 2444 6103 2451 6129
rect 2387 6102 2451 6103
rect 2174 6101 2509 6102
rect 2043 6099 2510 6101
rect 1731 6098 1779 6099
rect 2043 6098 2187 6099
rect 1731 6094 2187 6098
rect 2441 6097 2510 6099
rect 1731 6046 1745 6094
rect 1601 6033 1751 6046
rect 1601 5265 1608 6033
rect 2174 6046 2187 6094
rect 2174 6036 2175 6046
rect 2505 5902 2510 6097
rect 2574 5950 2581 6148
rect 2878 6145 2889 6148
rect 2600 6025 2635 6033
rect 2600 5968 2604 6025
rect 2580 5937 2581 5950
rect 2597 5903 2604 5968
rect 2880 5950 2887 6145
rect 3072 6085 3085 6153
rect 3245 6161 3276 6167
rect 3289 6161 3290 6172
rect 3449 6166 3450 6175
rect 3072 6074 3154 6085
rect 2906 6025 2941 6033
rect 2906 5968 2910 6025
rect 2886 5937 2887 5950
rect 2903 5903 2910 5968
rect 3072 5942 3085 6074
rect 3245 6085 3252 6161
rect 3186 6074 3252 6085
rect 3245 5963 3252 6074
rect 3271 6038 3306 6046
rect 3271 5981 3275 6038
rect 3251 5950 3252 5963
rect 3268 5916 3275 5981
rect 3437 5990 3450 6166
rect 3977 6110 3978 6119
rect 3977 6017 3989 6110
rect 4447 6116 4448 6125
rect 4447 6019 4459 6116
rect 4447 6018 4677 6019
rect 4265 6017 4677 6018
rect 3977 6016 4153 6017
rect 3977 6015 4217 6016
rect 3977 6012 4195 6015
rect 3795 6011 4195 6012
rect 3672 6009 3747 6010
rect 3672 6000 3725 6009
rect 3745 6000 3747 6009
rect 3815 6009 4195 6011
rect 3815 6000 3989 6009
rect 4142 6006 4195 6009
rect 4215 6006 4217 6015
rect 4285 6006 4677 6017
rect 4688 6006 4690 6019
rect 3437 5955 3450 5973
rect 3677 5949 3693 6000
rect 3266 5914 3275 5916
rect 3226 5909 3275 5914
rect 3226 5908 3285 5909
rect 2524 5902 2539 5903
rect 2505 5901 2539 5902
rect 2595 5901 2604 5903
rect 2505 5896 2604 5901
rect 2879 5901 2895 5902
rect 2901 5901 2910 5903
rect 2505 5895 2510 5896
rect 2527 5895 2614 5896
rect 2849 5896 2910 5901
rect 2849 5895 2920 5896
rect 2585 5868 2597 5895
rect 2879 5868 2895 5895
rect 3244 5868 3257 5908
rect 3677 5873 3692 5949
rect 3265 5868 3694 5873
rect 2585 5852 3694 5868
rect 3265 5851 3694 5852
rect 2894 5630 3845 5631
rect 2894 5626 3828 5630
rect 2893 5616 3828 5626
rect 2893 5391 2904 5616
rect 3977 5447 3978 5456
rect 3475 5401 3488 5404
rect 2901 5389 2904 5391
rect 3084 5392 3097 5395
rect 3292 5394 3314 5398
rect 2901 5386 2923 5389
rect 2559 5376 2581 5379
rect 2550 5368 2581 5376
rect 2594 5368 2595 5379
rect 2892 5378 2923 5386
rect 2936 5378 2937 5389
rect 3096 5383 3097 5392
rect 2043 5302 2050 5329
rect 2444 5306 2451 5338
rect 2169 5303 2451 5306
rect 2169 5302 2452 5303
rect 2043 5301 2452 5302
rect 1740 5298 2452 5301
rect 1740 5294 2174 5298
rect 1740 5265 1750 5294
rect 1783 5293 2050 5294
rect 2169 5287 2174 5294
rect 2167 5267 2175 5287
rect 1601 5261 1766 5265
rect 1601 5252 1752 5261
rect 2444 5123 2452 5298
rect 2550 5170 2557 5368
rect 2576 5245 2611 5253
rect 2576 5188 2580 5245
rect 2556 5157 2557 5170
rect 2573 5123 2580 5188
rect 2892 5180 2899 5378
rect 3084 5314 3097 5383
rect 3283 5387 3314 5394
rect 3327 5387 3328 5398
rect 3487 5392 3488 5401
rect 3084 5299 3186 5314
rect 3283 5314 3290 5387
rect 3221 5299 3290 5314
rect 2918 5255 2953 5263
rect 2918 5198 2922 5255
rect 2898 5167 2899 5180
rect 2915 5133 2922 5198
rect 3084 5172 3097 5299
rect 3283 5189 3290 5299
rect 3475 5274 3488 5392
rect 3977 5351 3989 5447
rect 4447 5453 4448 5462
rect 4447 5357 4459 5453
rect 4447 5355 4677 5357
rect 4265 5354 4677 5355
rect 4142 5352 4217 5353
rect 4142 5351 4195 5352
rect 3977 5349 4195 5351
rect 3795 5348 4195 5349
rect 3672 5346 3747 5347
rect 3672 5337 3725 5346
rect 3745 5337 3747 5346
rect 3815 5343 4195 5348
rect 4215 5343 4217 5352
rect 4285 5344 4677 5354
rect 4285 5343 4459 5344
rect 4688 5344 4690 5357
rect 3815 5337 3989 5343
rect 3681 5277 3698 5337
rect 3309 5264 3344 5272
rect 3309 5207 3313 5264
rect 3289 5176 3290 5189
rect 3306 5142 3313 5207
rect 3475 5181 3488 5257
rect 3682 5256 3698 5277
rect 3304 5140 3313 5142
rect 3265 5135 3313 5140
rect 3265 5134 3323 5135
rect 2913 5131 2922 5133
rect 2861 5126 2922 5131
rect 2861 5125 2932 5126
rect 2444 5121 2515 5123
rect 2571 5121 2580 5123
rect 2444 5116 2580 5121
rect 2444 5115 2590 5116
rect 2444 5114 2507 5115
rect 2560 5083 2569 5115
rect 2863 5083 2870 5125
rect 3282 5083 3293 5134
rect 3681 5084 3698 5256
rect 3314 5083 3700 5084
rect 2560 5069 3700 5083
rect 2863 5068 2870 5069
rect 3314 5064 3700 5069
<< m3contact >>
rect 3704 5583 3725 5605
<< m123contact >>
rect 2589 7890 2603 7900
rect 2687 7891 2699 7899
rect 3756 7997 3767 8015
rect 3222 7936 3233 7956
rect 3005 7896 3017 7904
rect 3323 7894 3335 7902
rect 2087 7797 2093 7802
rect 2653 7691 2660 7696
rect 2971 7696 2978 7701
rect 3289 7694 3296 7699
rect 3236 7645 3244 7659
rect 4026 7814 4039 7827
rect 4660 7814 4677 7826
rect 3722 7720 3742 7729
rect 3792 7720 3812 7731
rect 4192 7726 4212 7735
rect 4262 7726 4282 7737
rect 4669 7736 4690 7749
rect 2543 7520 2574 7535
rect 2712 7530 2719 7536
rect 3030 7535 3037 7541
rect 3348 7533 3355 7539
rect 4227 7644 4240 7660
rect 2542 7135 2575 7142
rect 2636 7136 2648 7144
rect 3758 7216 3771 7228
rect 3229 7190 3236 7198
rect 2990 7151 3002 7159
rect 3333 7149 3345 7157
rect 2082 7040 2091 7045
rect 2602 6936 2609 6941
rect 3162 6979 3191 6993
rect 2956 6951 2963 6956
rect 3299 6949 3306 6954
rect 4035 7021 4046 7036
rect 4680 7022 4691 7036
rect 3439 6895 3451 6911
rect 3725 6948 3745 6957
rect 3795 6948 3815 6959
rect 4195 6954 4215 6963
rect 4265 6954 4285 6965
rect 4677 6955 4688 6970
rect 2661 6775 2668 6781
rect 3015 6790 3022 6796
rect 3358 6788 3365 6794
rect 2528 6672 2547 6689
rect 2547 6236 2574 6254
rect 2660 6245 2672 6253
rect 3709 6342 3731 6364
rect 3226 6303 3241 6318
rect 3331 6258 3343 6266
rect 2966 6245 2978 6253
rect 2086 6150 2094 6155
rect 2626 6045 2633 6050
rect 2932 6045 2939 6050
rect 3154 6072 3186 6086
rect 3297 6058 3304 6063
rect 4027 6071 4037 6085
rect 4672 6071 4683 6084
rect 3725 6000 3745 6009
rect 3795 6000 3815 6011
rect 4195 6006 4215 6015
rect 4265 6006 4285 6017
rect 4677 6005 4688 6020
rect 3437 5973 3451 5990
rect 2531 5860 2557 5875
rect 2685 5884 2692 5890
rect 2991 5884 2998 5890
rect 3356 5897 3363 5903
rect 2530 5458 2556 5473
rect 2636 5465 2648 5473
rect 3262 5535 3286 5560
rect 3369 5484 3381 5492
rect 2978 5475 2990 5483
rect 2087 5370 2094 5375
rect 2602 5265 2609 5270
rect 3186 5299 3221 5315
rect 2944 5275 2951 5280
rect 3335 5284 3342 5289
rect 4031 5416 4037 5429
rect 4668 5414 4686 5428
rect 3725 5337 3745 5346
rect 3795 5337 3815 5348
rect 4195 5343 4215 5352
rect 4265 5343 4285 5354
rect 4677 5343 4688 5358
rect 3475 5257 3489 5274
rect 2661 5104 2668 5110
rect 3003 5114 3010 5120
rect 3394 5123 3401 5129
<< metal3 >>
rect 3750 8021 3778 8023
rect 2831 8015 3778 8021
rect 2831 7997 3756 8015
rect 3767 7997 3778 8015
rect 2833 7988 2854 7997
rect 3750 7996 3778 7997
rect 2834 7959 2854 7988
rect 2278 7951 2319 7953
rect 2833 7951 2854 7959
rect 2086 7929 2913 7951
rect 3221 7936 3222 7956
rect 2088 7881 2095 7929
rect 2278 7928 2319 7929
rect 2902 7904 2911 7929
rect 2087 7802 2095 7881
rect 2093 7799 2095 7802
rect 2583 7890 2589 7899
rect 2603 7891 2687 7899
rect 2603 7890 2699 7891
rect 2901 7896 3005 7904
rect 3221 7902 3233 7936
rect 2901 7895 3017 7896
rect 2901 7894 2911 7895
rect 3219 7894 3323 7902
rect 2087 7795 2093 7797
rect 2583 7760 2590 7890
rect 2901 7765 2908 7894
rect 2582 7752 2590 7760
rect 2888 7757 2908 7765
rect 3219 7893 3335 7894
rect 3219 7892 3233 7893
rect 3219 7763 3226 7892
rect 4039 7814 4660 7826
rect 4026 7813 4677 7814
rect 2583 7695 2590 7752
rect 2901 7700 2908 7757
rect 3218 7755 3226 7763
rect 2901 7696 2971 7700
rect 3219 7698 3226 7755
rect 2583 7691 2653 7695
rect 2583 7536 2590 7691
rect 2901 7541 2908 7696
rect 3219 7694 3289 7698
rect 2543 7535 2712 7536
rect 2574 7530 2712 7535
rect 2901 7535 3030 7541
rect 3219 7539 3226 7694
rect 3235 7645 3236 7659
rect 3244 7645 4227 7659
rect 4240 7645 4260 7659
rect 2901 7534 2908 7535
rect 3219 7533 3348 7539
rect 3219 7532 3226 7533
rect 2574 7527 2595 7530
rect 2574 7520 2591 7527
rect 2885 7224 3758 7228
rect 2884 7216 3758 7224
rect 3771 7216 3772 7228
rect 2884 7215 3772 7216
rect 2884 7163 2898 7215
rect 2080 7159 2898 7163
rect 3229 7198 3237 7199
rect 3236 7190 3237 7198
rect 2080 7151 2990 7159
rect 2080 7150 2560 7151
rect 2574 7150 3002 7151
rect 3229 7157 3237 7190
rect 2082 7119 2093 7150
rect 2081 7103 2093 7119
rect 2532 7143 2560 7144
rect 2574 7143 2636 7144
rect 2532 7142 2636 7143
rect 2532 7135 2542 7142
rect 2575 7136 2636 7142
rect 2575 7135 2648 7136
rect 2532 7123 2540 7135
rect 2081 7045 2091 7103
rect 2081 7042 2082 7045
rect 2082 7008 2091 7040
rect 2532 7005 2539 7123
rect 2886 7020 2893 7150
rect 3229 7149 3333 7157
rect 3229 7148 3345 7149
rect 3229 7146 3237 7148
rect 3229 7068 3236 7146
rect 3230 7058 3236 7068
rect 2873 7012 2893 7020
rect 2528 6997 2539 7005
rect 2532 6940 2539 6997
rect 2886 6955 2893 7012
rect 2886 6951 2956 6955
rect 3229 6953 3236 7058
rect 4034 7022 4035 7036
rect 4046 7022 4680 7036
rect 2532 6936 2602 6940
rect 2532 6782 2539 6936
rect 2886 6796 2893 6951
rect 3229 6949 3299 6953
rect 2886 6790 3015 6796
rect 3229 6794 3236 6949
rect 3439 6911 3456 6913
rect 3451 6897 3456 6911
rect 2886 6789 2893 6790
rect 3229 6788 3358 6794
rect 3229 6787 3236 6788
rect 2532 6781 2554 6782
rect 2532 6776 2661 6781
rect 2527 6775 2661 6776
rect 2527 6772 2554 6775
rect 2527 6689 2546 6772
rect 2527 6673 2528 6689
rect 2883 6364 2899 6370
rect 2883 6343 3709 6364
rect 2528 6274 2576 6275
rect 2883 6274 2899 6343
rect 3731 6343 3732 6364
rect 3227 6318 3244 6319
rect 3241 6303 3244 6318
rect 2086 6270 2904 6274
rect 2086 6261 2907 6270
rect 2088 6231 2099 6261
rect 2574 6253 2580 6254
rect 2860 6253 2907 6261
rect 3227 6266 3244 6303
rect 3227 6258 3331 6266
rect 3227 6257 3343 6258
rect 2574 6245 2660 6253
rect 2860 6251 2966 6253
rect 2574 6244 2672 6245
rect 2862 6245 2966 6251
rect 2862 6244 2978 6245
rect 3227 6252 3244 6257
rect 2087 6219 2099 6231
rect 2556 6235 2567 6236
rect 2556 6228 2565 6235
rect 2087 6155 2096 6219
rect 2094 6153 2096 6155
rect 2086 6117 2094 6150
rect 2556 6114 2563 6228
rect 2862 6114 2869 6244
rect 3227 6195 3234 6252
rect 3226 6178 3234 6195
rect 3226 6167 3233 6178
rect 3226 6160 3234 6167
rect 3227 6127 3234 6160
rect 3226 6119 3234 6127
rect 2547 6106 2563 6114
rect 2849 6106 2869 6114
rect 2556 6049 2563 6106
rect 2556 6045 2626 6049
rect 2862 6049 2869 6106
rect 3227 6062 3234 6119
rect 4037 6071 4672 6084
rect 4683 6071 4684 6084
rect 4027 6070 4684 6071
rect 3227 6058 3297 6062
rect 2862 6045 2932 6049
rect 2556 5915 2563 6045
rect 2556 5894 2564 5915
rect 2518 5890 2575 5894
rect 2862 5890 2869 6045
rect 3227 5903 3234 6058
rect 3437 5990 3485 5991
rect 3451 5973 3485 5990
rect 3227 5897 3356 5903
rect 3227 5896 3234 5897
rect 2518 5884 2685 5890
rect 2862 5884 2991 5890
rect 2518 5875 2575 5884
rect 2862 5883 2869 5884
rect 2518 5860 2531 5875
rect 2557 5860 2575 5875
rect 2870 5584 3704 5605
rect 2087 5490 2098 5491
rect 2871 5490 2881 5584
rect 3262 5560 3282 5561
rect 3262 5492 3282 5535
rect 2085 5489 2533 5490
rect 2551 5489 2903 5490
rect 2085 5483 2903 5489
rect 3262 5484 3369 5492
rect 3262 5483 3381 5484
rect 2085 5478 2978 5483
rect 2085 5477 2533 5478
rect 2551 5477 2978 5478
rect 2087 5438 2098 5477
rect 2874 5475 2978 5477
rect 3262 5477 3282 5483
rect 2874 5474 2990 5475
rect 2556 5465 2636 5473
rect 2556 5464 2648 5465
rect 2556 5458 2557 5464
rect 2087 5375 2096 5438
rect 2094 5370 2096 5375
rect 2087 5368 2096 5370
rect 2532 5334 2539 5458
rect 2874 5344 2881 5474
rect 2861 5336 2881 5344
rect 2529 5323 2539 5334
rect 2532 5269 2539 5323
rect 2874 5279 2881 5336
rect 3265 5288 3272 5477
rect 4030 5416 4031 5429
rect 4037 5428 4687 5429
rect 4037 5416 4668 5428
rect 4030 5415 4668 5416
rect 4686 5415 4687 5428
rect 3265 5284 3335 5288
rect 2874 5275 2944 5279
rect 2532 5265 2602 5269
rect 2532 5110 2539 5265
rect 2874 5120 2881 5275
rect 3265 5129 3272 5284
rect 3489 5257 3492 5274
rect 3265 5123 3394 5129
rect 3265 5122 3272 5123
rect 2874 5114 3003 5120
rect 2874 5113 2881 5114
rect 2532 5104 2661 5110
rect 2532 5103 2539 5104
<< labels >>
rlabel metal1 1669 7840 1669 7840 1 vdd
rlabel metal2 1606 7681 1606 7681 1 gnd
rlabel metal1 2800 5385 2800 5385 1 bs3
rlabel metal1 2781 6101 2781 6101 1 bs2
rlabel metal1 2763 7006 2763 7006 1 bs1
rlabel metal1 2800 7737 2800 7737 1 bs0
rlabel metal2 3156 7746 3156 7746 1 axorb
rlabel polysilicon 1691 8332 1708 8345 1 D1
rlabel polysilicon 1782 8332 1799 8345 1 D0
rlabel metal1 3386 7803 3441 7810 1 OUT_AS0
rlabel metal1 3396 7058 3451 7065 1 OUT_AS1
rlabel metal1 3394 6167 3449 6174 1 OUT_AS2
rlabel metal1 4980 5419 4988 5422 1 C
rlabel polysilicon 1821 7761 1829 7767 1 ASA0
rlabel polysilicon 2106 7865 2117 7872 1 DAS
rlabel polysilicon 1819 7015 1828 7021 1 ASA1
rlabel polysilicon 1820 6109 1829 6115 1 ASA2
rlabel polysilicon 1818 5328 1827 5334 1 ASA3
rlabel polysilicon 2220 5334 2228 5338 1 ASB3
rlabel polysilicon 2221 6122 2229 6126 1 ASB2
rlabel polysilicon 2221 7006 2229 7010 1 ASB1
rlabel polysilicon 2218 7762 2226 7766 1 ASB0
rlabel metal1 3433 5393 3475 5400 1 OUT_AS3
<< end >>
