magic
tech scmos
timestamp 1701790942
<< nwell >>
rect 767 384 803 416
rect 767 338 803 370
rect 855 331 891 363
rect 343 229 379 261
rect 399 229 435 261
rect 454 220 490 252
rect 560 229 596 261
rect 616 229 652 261
rect 671 220 707 252
rect 307 58 329 86
rect 425 83 447 111
rect 377 54 399 82
rect 562 60 584 88
rect 680 85 702 113
rect 632 56 654 84
rect 448 4 470 32
rect 703 6 725 34
<< ntransistor >>
rect 386 183 390 203
rect 773 298 777 318
rect 824 298 828 318
rect 871 301 875 321
rect 470 190 474 210
rect 386 143 390 163
rect 603 183 607 203
rect 687 190 691 210
rect 603 143 607 163
rect 454 95 464 99
rect 709 97 719 101
rect 313 39 323 43
rect 383 35 393 39
rect 431 16 441 20
rect 568 41 578 45
rect 638 37 648 41
rect 686 18 696 22
<< ptransistor >>
rect 784 390 786 410
rect 360 235 362 255
rect 416 235 418 255
rect 471 226 473 246
rect 784 344 786 364
rect 872 337 874 357
rect 577 235 579 255
rect 633 235 635 255
rect 688 226 690 246
rect 431 96 441 98
rect 686 98 696 100
rect 313 71 323 73
rect 383 67 393 69
rect 568 73 578 75
rect 638 69 648 71
rect 454 17 464 19
rect 709 19 719 21
<< ndiffusion >>
rect 385 183 386 203
rect 390 183 391 203
rect 772 298 773 318
rect 777 298 778 318
rect 823 298 824 318
rect 828 298 829 318
rect 870 301 871 321
rect 875 301 876 321
rect 469 190 470 210
rect 474 190 475 210
rect 385 143 386 163
rect 390 143 391 163
rect 454 99 464 100
rect 602 183 603 203
rect 607 183 608 203
rect 686 190 687 210
rect 691 190 692 210
rect 602 143 603 163
rect 607 143 608 163
rect 709 101 719 102
rect 454 94 464 95
rect 709 96 719 97
rect 313 43 323 44
rect 383 39 393 40
rect 313 38 323 39
rect 383 34 393 35
rect 431 20 441 21
rect 431 15 441 16
rect 568 45 578 46
rect 638 41 648 42
rect 568 40 578 41
rect 638 36 648 37
rect 686 22 696 23
rect 686 17 696 18
<< pdiffusion >>
rect 783 390 784 410
rect 786 390 787 410
rect 359 235 360 255
rect 362 235 363 255
rect 415 235 416 255
rect 418 235 419 255
rect 470 226 471 246
rect 473 226 474 246
rect 783 344 784 364
rect 786 344 787 364
rect 871 337 872 357
rect 874 337 875 357
rect 576 235 577 255
rect 579 235 580 255
rect 632 235 633 255
rect 635 235 636 255
rect 687 226 688 246
rect 690 226 691 246
rect 431 98 441 100
rect 431 94 441 96
rect 686 100 696 102
rect 313 73 323 75
rect 313 69 323 71
rect 383 69 393 71
rect 383 65 393 67
rect 686 96 696 98
rect 568 75 578 77
rect 568 71 578 73
rect 638 71 648 73
rect 638 67 648 69
rect 454 19 464 21
rect 454 15 464 17
rect 709 21 719 23
rect 709 17 719 19
<< ndcontact >>
rect 375 183 385 203
rect 391 183 401 203
rect 762 298 772 318
rect 778 298 788 318
rect 813 298 823 318
rect 829 298 839 318
rect 860 301 870 321
rect 876 301 886 321
rect 459 190 469 210
rect 475 190 485 210
rect 375 143 385 163
rect 391 143 401 163
rect 454 100 464 105
rect 592 183 602 203
rect 608 183 618 203
rect 676 190 686 210
rect 692 190 702 210
rect 592 143 602 163
rect 608 143 618 163
rect 709 102 719 107
rect 454 89 464 94
rect 709 91 719 96
rect 313 44 323 49
rect 383 40 393 45
rect 313 33 323 38
rect 383 29 393 34
rect 431 21 441 26
rect 431 10 441 15
rect 568 46 578 51
rect 638 42 648 47
rect 568 35 578 40
rect 638 31 648 36
rect 686 23 696 28
rect 686 12 696 17
<< pdcontact >>
rect 773 390 783 410
rect 787 390 797 410
rect 349 235 359 255
rect 363 235 373 255
rect 405 235 415 255
rect 419 235 429 255
rect 460 226 470 246
rect 474 226 484 246
rect 773 344 783 364
rect 787 344 797 364
rect 861 337 871 357
rect 875 337 885 357
rect 566 235 576 255
rect 580 235 590 255
rect 622 235 632 255
rect 636 235 646 255
rect 677 226 687 246
rect 691 226 701 246
rect 431 100 441 105
rect 686 102 696 107
rect 431 89 441 94
rect 313 75 323 80
rect 383 71 393 76
rect 313 64 323 69
rect 383 60 393 65
rect 686 91 696 96
rect 568 77 578 82
rect 638 73 648 78
rect 568 66 578 71
rect 638 62 648 67
rect 454 21 464 26
rect 454 10 464 15
rect 709 23 719 28
rect 709 12 719 17
<< psubstratepcontact >>
rect 742 284 746 288
rect 835 284 839 288
rect 855 284 859 288
rect 887 284 891 288
rect 343 133 347 137
rect 431 133 435 137
rect 454 133 458 137
rect 486 133 490 137
rect 560 133 564 137
rect 648 133 652 137
rect 671 133 675 137
rect 703 133 707 137
rect 316 25 320 29
rect 386 21 390 25
rect 571 27 575 31
rect 641 23 645 27
<< nsubstratencontact >>
rect 767 416 771 420
rect 799 416 803 420
rect 855 416 859 420
rect 887 416 891 420
rect 343 261 347 265
rect 431 261 435 265
rect 454 261 458 265
rect 486 261 490 265
rect 560 261 564 265
rect 648 261 652 265
rect 671 261 675 265
rect 703 261 707 265
rect 434 111 438 115
rect 689 113 693 117
rect 316 86 320 90
rect 386 82 390 86
rect 571 88 575 92
rect 641 84 645 88
rect 457 32 461 36
rect 712 34 716 38
<< polysilicon >>
rect 784 410 786 413
rect 784 381 786 390
rect 494 377 735 381
rect 771 377 786 381
rect 360 255 362 258
rect 416 255 418 258
rect 471 246 473 249
rect 360 226 362 235
rect 416 226 418 235
rect 347 222 362 226
rect 403 222 418 226
rect 375 206 390 210
rect 386 203 390 206
rect 386 180 390 183
rect 414 170 418 222
rect 471 217 473 226
rect 456 215 473 217
rect 494 217 498 377
rect 784 364 786 367
rect 872 357 874 360
rect 784 335 786 344
rect 771 331 811 335
rect 773 318 777 321
rect 773 295 777 298
rect 760 291 777 295
rect 807 295 811 331
rect 872 328 874 337
rect 857 326 874 328
rect 857 324 875 326
rect 871 321 875 324
rect 824 318 828 321
rect 871 298 875 301
rect 824 295 828 298
rect 807 291 828 295
rect 577 255 579 258
rect 633 255 635 258
rect 688 246 690 249
rect 577 226 579 235
rect 633 226 635 235
rect 564 222 579 226
rect 620 222 635 226
rect 456 213 474 215
rect 470 210 474 213
rect 592 206 607 210
rect 470 187 474 190
rect 375 166 418 170
rect 386 163 390 166
rect 386 140 390 143
rect 545 101 550 206
rect 603 203 607 206
rect 603 180 607 183
rect 631 170 635 222
rect 688 217 690 226
rect 673 215 690 217
rect 673 213 691 215
rect 687 210 691 213
rect 687 187 691 190
rect 592 166 635 170
rect 603 163 607 166
rect 603 140 607 143
rect 342 96 431 98
rect 441 96 444 98
rect 451 95 454 99
rect 464 98 467 99
rect 464 96 476 98
rect 597 98 686 100
rect 696 98 699 100
rect 464 95 467 96
rect 329 86 347 90
rect 343 82 377 86
rect 305 71 313 73
rect 323 71 326 73
rect 375 67 383 69
rect 393 67 396 69
rect 474 57 476 96
rect 706 97 709 101
rect 719 100 722 101
rect 719 98 731 100
rect 719 97 722 98
rect 584 88 602 92
rect 598 84 632 88
rect 560 73 568 75
rect 578 73 581 75
rect 630 69 638 71
rect 648 69 651 71
rect 729 59 731 98
rect 729 57 739 59
rect 474 55 484 57
rect 310 42 313 43
rect 305 40 313 42
rect 310 39 313 40
rect 323 39 326 43
rect 380 38 383 39
rect 375 36 383 38
rect 380 35 383 36
rect 393 35 396 39
rect 328 25 364 29
rect 428 18 431 20
rect 342 16 431 18
rect 441 16 444 20
rect 474 19 476 55
rect 451 17 454 19
rect 464 17 476 19
rect 482 3 484 55
rect 565 44 568 45
rect 560 42 568 44
rect 565 41 568 42
rect 578 41 581 45
rect 635 40 638 41
rect 630 38 638 40
rect 635 37 638 38
rect 648 37 651 41
rect 583 27 619 31
rect 683 20 686 22
rect 597 18 686 20
rect 696 18 699 22
rect 729 21 731 57
rect 706 19 709 21
rect 719 19 731 21
rect 349 1 484 3
rect 737 5 739 57
rect 604 3 739 5
<< polycontact >>
rect 735 377 739 381
rect 767 377 771 381
rect 343 222 347 226
rect 371 206 375 210
rect 452 213 456 217
rect 767 331 771 335
rect 756 291 760 295
rect 853 324 857 328
rect 560 222 564 226
rect 494 213 498 217
rect 545 206 550 210
rect 588 206 592 210
rect 371 166 375 170
rect 338 95 342 99
rect 669 213 673 217
rect 588 166 592 170
rect 545 97 550 101
rect 593 97 597 101
rect 325 86 329 90
rect 377 82 381 86
rect 301 70 305 74
rect 371 66 375 70
rect 580 88 584 92
rect 632 84 636 88
rect 556 72 560 76
rect 626 68 630 72
rect 301 39 305 43
rect 371 35 375 39
rect 323 25 328 29
rect 364 25 369 29
rect 338 15 342 19
rect 345 0 349 4
rect 556 41 560 45
rect 626 37 630 41
rect 578 27 583 31
rect 619 27 624 31
rect 593 17 597 21
rect 600 2 604 6
<< metal1 >>
rect 699 416 767 420
rect 771 416 799 420
rect 803 416 855 420
rect 859 416 887 420
rect 699 265 703 416
rect 773 410 783 416
rect 739 377 767 381
rect 735 335 739 377
rect 787 374 797 390
rect 767 370 803 374
rect 773 364 783 370
rect 715 331 767 335
rect 347 261 431 265
rect 435 261 438 265
rect 349 255 359 261
rect 405 255 415 261
rect 444 261 454 265
rect 458 261 486 265
rect 490 261 560 265
rect 564 261 648 265
rect 652 261 671 265
rect 675 261 703 265
rect 276 222 343 226
rect 276 56 281 222
rect 328 210 332 222
rect 363 217 373 235
rect 419 217 429 235
rect 460 246 470 261
rect 566 255 576 261
rect 622 255 632 261
rect 475 217 484 226
rect 545 222 560 226
rect 343 213 452 217
rect 475 213 494 217
rect 328 206 371 210
rect 391 203 401 213
rect 475 210 484 213
rect 545 210 550 222
rect 580 217 590 235
rect 636 217 646 235
rect 677 246 687 261
rect 692 217 701 226
rect 715 217 719 331
rect 735 295 739 331
rect 787 328 797 344
rect 861 357 871 416
rect 876 328 885 337
rect 742 324 853 328
rect 876 324 899 328
rect 762 318 772 324
rect 813 318 823 324
rect 876 321 885 324
rect 735 291 756 295
rect 778 288 788 298
rect 829 288 839 298
rect 860 288 870 301
rect 560 213 669 217
rect 692 213 719 217
rect 735 284 742 288
rect 746 284 835 288
rect 839 284 855 288
rect 859 284 887 288
rect 550 206 588 210
rect 608 203 618 213
rect 692 210 701 213
rect 375 177 385 183
rect 375 173 401 177
rect 358 166 371 170
rect 391 163 401 173
rect 375 137 385 143
rect 459 137 469 190
rect 592 177 602 183
rect 592 173 618 177
rect 578 166 588 170
rect 608 163 618 173
rect 592 137 602 143
rect 676 137 686 190
rect 735 137 739 284
rect 347 133 431 137
rect 435 133 454 137
rect 458 133 486 137
rect 490 133 560 137
rect 564 133 648 137
rect 652 133 671 137
rect 675 133 703 137
rect 707 133 739 137
rect 429 115 447 116
rect 429 111 434 115
rect 438 111 447 115
rect 684 117 697 118
rect 684 113 689 117
rect 693 113 697 117
rect 441 100 454 105
rect 464 100 502 105
rect 696 102 709 107
rect 719 102 757 107
rect 286 95 338 99
rect 286 56 290 95
rect 307 86 316 90
rect 320 86 325 90
rect 363 89 431 94
rect 441 89 454 94
rect 316 80 320 86
rect 301 56 305 70
rect 276 52 305 56
rect 286 19 290 52
rect 301 43 305 52
rect 316 56 320 64
rect 316 52 349 56
rect 363 56 367 89
rect 381 82 386 86
rect 390 82 410 86
rect 386 76 390 82
rect 411 76 416 81
rect 411 70 453 76
rect 371 56 375 66
rect 363 52 375 56
rect 316 49 320 52
rect 316 29 320 33
rect 313 25 316 29
rect 320 25 323 29
rect 286 15 338 19
rect 345 4 349 52
rect 371 39 375 52
rect 386 52 390 60
rect 386 48 411 52
rect 386 45 390 48
rect 386 25 390 29
rect 407 26 411 48
rect 448 36 453 70
rect 498 58 502 100
rect 541 58 545 101
rect 550 97 593 101
rect 562 88 571 92
rect 575 88 580 92
rect 618 91 686 96
rect 696 91 709 96
rect 571 82 575 88
rect 556 58 560 72
rect 498 54 560 58
rect 448 32 457 36
rect 461 32 470 36
rect 364 21 386 25
rect 390 21 393 25
rect 407 21 431 26
rect 441 21 454 26
rect 386 -6 390 21
rect 498 15 502 54
rect 541 21 545 54
rect 556 45 560 54
rect 571 58 575 66
rect 571 54 604 58
rect 618 58 622 91
rect 636 84 641 88
rect 645 84 665 88
rect 641 78 645 84
rect 666 78 671 83
rect 666 72 708 78
rect 626 58 630 68
rect 618 54 630 58
rect 571 51 575 54
rect 571 31 575 35
rect 568 27 571 31
rect 575 27 578 31
rect 541 17 593 21
rect 441 10 454 15
rect 464 10 502 15
rect 600 6 604 54
rect 626 41 630 54
rect 641 54 645 62
rect 641 50 666 54
rect 641 47 645 50
rect 641 27 645 31
rect 662 28 666 50
rect 703 38 708 72
rect 753 60 757 102
rect 753 54 766 60
rect 703 34 712 38
rect 716 34 725 38
rect 619 23 641 27
rect 645 23 648 27
rect 662 23 686 28
rect 696 23 709 28
rect 621 -6 625 23
rect 753 17 757 54
rect 696 12 709 17
rect 719 12 757 17
rect 789 -6 793 284
rect 386 -10 865 -6
<< m2contact >>
rect 353 166 358 171
rect 423 111 429 116
rect 678 113 684 118
rect 358 52 363 57
rect 410 81 416 86
rect 613 54 618 59
rect 665 83 671 88
<< metal2 >>
rect 353 52 358 166
rect 573 119 578 165
rect 416 111 423 116
rect 573 114 614 119
rect 410 86 416 111
rect 609 59 614 114
rect 665 113 678 118
rect 665 88 671 113
rect 609 54 613 59
<< m123contact >>
rect 438 259 444 265
rect 573 165 578 170
rect 410 111 416 116
rect 697 113 702 118
<< metal3 >>
rect 438 143 444 259
rect 535 165 573 170
rect 410 138 444 143
rect 410 129 416 138
rect 410 125 702 129
rect 410 116 416 125
rect 697 118 702 125
<< labels >>
rlabel metal1 328 222 347 226 1 A
rlabel metal1 757 54 766 60 7 S1
rlabel metal3 535 165 545 170 1 Cin
rlabel metal1 343 133 707 137 1 Gnd
rlabel metal1 343 261 707 265 5 VDD
rlabel metal1 885 324 899 328 1 C
rlabel metal1 356 166 375 170 1 B
<< end >>
