* SPICE3 file created from OUTble.ext - technology: scmos

.include TSMC_180nm.txt
.param SUPPLY = 1.8
.global Gnd
Vdd VDD Gnd 'SUPPLY'
.option scale=0.09u

VinIn1 In1 Gnd DC 'SUPPLY'
VinIn2 In2 Gnd DC 'SUPPLY'
VinIn3 In3 Gnd DC 'SUPPLY'
VinIn4 In4 Gnd DC 'SUPPLY'
VinIn5 In5 Gnd DC 'SUPPLY'
VinIn6 In6 Gnd DC 'SUPPLY'
VinIn7 In7 Gnd DC 0
VinIn8 In8 Gnd DC 0

VinD1 EN Gnd PULSE('SUPPLY' 0 0ns 100ps 100ps 5n 10n)

M1000 a_964_407# EN VDD VDD CMOSP w=20 l=2
+  ad=440 pd=124 as=5280 ps=1488
M1001 a_1561_407# In5 VDD VDD CMOSP w=20 l=2
+  ad=440 pd=124 as=0 ps=0
M1002 OUT7 a_1968_407# VDD w_2060_392# CMOSP w=20 l=2
+  ad=220 pd=62 as=0 ps=0
M1003 OUT8 a_2171_407# VDD w_2263_392# CMOSP w=20 l=2
+  ad=220 pd=62 as=0 ps=0
M1004 a_1561_407# EN VDD VDD CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1005 a_1764_407# EN VDD VDD CMOSP w=20 l=2
+  ad=440 pd=124 as=0 ps=0
M1006 a_1968_407# EN a_1981_355# Gnd CMOSN w=20 l=4
+  ad=220 pd=62 as=440 ps=124
M1007 a_1169_355# In3 Gnd Gnd CMOSN w=20 l=4
+  ad=440 pd=124 as=3520 ps=992
M1008 a_1371_355# In4 Gnd Gnd CMOSN w=20 l=4
+  ad=440 pd=124 as=0 ps=0
M1009 OUT8 a_2171_407# Gnd Gnd CMOSN w=20 l=4
+  ad=220 pd=62 as=0 ps=0
M1010 OUT1 a_766_407# VDD w_858_392# CMOSP w=20 l=2
+  ad=220 pd=62 as=0 ps=0
M1011 OUT2 a_964_407# VDD w_1056_392# CMOSP w=20 l=2
+  ad=220 pd=62 as=0 ps=0
M1012 a_2171_407# EN a_2184_355# Gnd CMOSN w=20 l=4
+  ad=220 pd=62 as=440 ps=124
M1013 OUT6 a_1764_407# VDD w_1856_392# CMOSP w=20 l=2
+  ad=220 pd=62 as=0 ps=0
M1014 a_1156_407# In3 VDD VDD CMOSP w=20 l=2
+  ad=440 pd=124 as=0 ps=0
M1015 a_1358_407# In4 VDD VDD CMOSP w=20 l=2
+  ad=440 pd=124 as=0 ps=0
M1016 a_1156_407# EN VDD VDD CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1017 a_1358_407# EN VDD VDD CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1018 a_964_407# EN a_977_355# Gnd CMOSN w=20 l=4
+  ad=220 pd=62 as=440 ps=124
M1019 a_1764_407# EN a_1777_355# Gnd CMOSN w=20 l=4
+  ad=220 pd=62 as=440 ps=124
M1020 a_1981_355# In7 Gnd Gnd CMOSN w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1021 OUT7 a_1968_407# Gnd Gnd CMOSN w=20 l=4
+  ad=220 pd=62 as=0 ps=0
M1022 a_2184_355# In8 Gnd Gnd CMOSN w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1023 OUT3 a_1156_407# VDD w_1248_392# CMOSP w=20 l=2
+  ad=220 pd=62 as=0 ps=0
M1024 OUT4 a_1358_407# VDD w_1450_392# CMOSP w=20 l=2
+  ad=220 pd=62 as=0 ps=0
M1025 OUT5 a_1561_407# VDD w_1653_392# CMOSP w=20 l=2
+  ad=220 pd=62 as=0 ps=0
M1026 OUT1 a_766_407# Gnd Gnd CMOSN w=20 l=4
+  ad=220 pd=62 as=0 ps=0
M1027 OUT2 a_964_407# Gnd Gnd CMOSN w=20 l=4
+  ad=220 pd=62 as=0 ps=0
M1028 a_1968_407# EN VDD VDD CMOSP w=20 l=2
+  ad=440 pd=124 as=0 ps=0
M1029 OUT5 a_1561_407# Gnd Gnd CMOSN w=20 l=4
+  ad=220 pd=62 as=0 ps=0
M1030 a_766_407# EN a_779_355# Gnd CMOSN w=20 l=4
+  ad=220 pd=62 as=440 ps=124
M1031 OUT6 a_1764_407# Gnd Gnd CMOSN w=20 l=4
+  ad=220 pd=62 as=0 ps=0
M1032 a_977_355# In2 Gnd Gnd CMOSN w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1033 a_2171_407# In8 VDD VDD CMOSP w=20 l=2
+  ad=440 pd=124 as=0 ps=0
M1034 a_1561_407# EN a_1574_355# Gnd CMOSN w=20 l=4
+  ad=220 pd=62 as=440 ps=124
M1035 a_1777_355# In6 Gnd Gnd CMOSN w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1036 a_2171_407# EN VDD VDD CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1037 a_964_407# In2 VDD VDD CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1038 a_1764_407# In6 VDD VDD CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1039 a_779_355# In1 Gnd Gnd CMOSN w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1040 OUT3 a_1156_407# Gnd Gnd CMOSN w=20 l=4
+  ad=220 pd=62 as=0 ps=0
M1041 OUT4 a_1358_407# Gnd Gnd CMOSN w=20 l=4
+  ad=220 pd=62 as=0 ps=0
M1042 a_1156_407# EN a_1169_355# Gnd CMOSN w=20 l=4
+  ad=220 pd=62 as=0 ps=0
M1043 a_1358_407# EN a_1371_355# Gnd CMOSN w=20 l=4
+  ad=220 pd=62 as=0 ps=0
M1044 a_1574_355# In5 Gnd Gnd CMOSN w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1045 a_1968_407# In7 VDD VDD CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1046 a_766_407# In1 VDD VDD CMOSP w=20 l=2
+  ad=440 pd=124 as=0 ps=0
M1047 a_766_407# EN VDD VDD CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
C0 VDD a_2171_407# 0.67fF
C1 EN a_1561_407# 0.47fF
C2 w_1856_392# a_1764_407# 0.06fF
C3 EN a_1358_407# 0.47fF
C4 w_1653_392# OUT5 0.06fF
C5 VDD a_1968_407# 0.67fF
C6 In5 a_1574_355# 0.19fF
C7 EN a_1156_407# 0.47fF
C8 VDD a_1764_407# 0.67fF
C9 a_1358_407# a_1371_355# 0.21fF
C10 EN a_766_407# 0.47fF
C11 VDD a_1561_407# 0.67fF
C12 EN a_964_407# 0.47fF
C13 VDD a_1358_407# 0.67fF
C14 w_1248_392# a_1156_407# 0.06fF
C15 VDD a_1156_407# 0.67fF
C16 w_1056_392# OUT2 0.06fF
C17 In2 a_977_355# 0.19fF
C18 OUT1 Gnd 0.14fF
C19 VDD a_766_407# 0.67fF
C20 Gnd a_1777_355# 0.21fF
C21 VDD a_964_407# 0.67fF
C22 VDD OUT1 0.21fF
C23 VDD w_2263_392# 0.06fF
C24 w_2263_392# a_2171_407# 0.06fF
C25 Gnd a_1169_355# 0.21fF
C26 VDD w_1653_392# 0.06fF
C27 w_2060_392# OUT7 0.06fF
C28 a_779_355# Gnd 0.21fF
C29 In7 a_1981_355# 0.19fF
C30 VDD w_1056_392# 0.06fF
C31 a_1764_407# a_1777_355# 0.21fF
C32 VDD In8 0.06fF
C33 In8 a_2171_407# 0.10fF
C34 w_1653_392# a_1561_407# 0.06fF
C35 VDD In7 0.06fF
C36 VDD In6 0.06fF
C37 w_1450_392# OUT4 0.06fF
C38 In4 a_1371_355# 0.19fF
C39 In7 a_1968_407# 0.10fF
C40 VDD In5 0.06fF
C41 a_1156_407# a_1169_355# 0.21fF
C42 VDD In4 0.06fF
C43 In6 a_1764_407# 0.10fF
C44 a_766_407# a_779_355# 0.21fF
C45 Gnd a_2184_355# 0.21fF
C46 VDD In3 0.06fF
C47 w_1056_392# a_964_407# 0.06fF
C48 VDD In1 0.06fF
C49 a_2171_407# a_2184_355# 0.21fF
C50 Gnd a_1574_355# 0.21fF
C51 VDD In2 0.06fF
C52 In5 a_1561_407# 0.10fF
C53 VDD w_2060_392# 0.06fF
C54 Gnd a_977_355# 0.21fF
C55 VDD w_1450_392# 0.06fF
C56 w_2060_392# a_1968_407# 0.06fF
C57 OUT8 Gnd 0.14fF
C58 In4 a_1358_407# 0.10fF
C59 VDD w_858_392# 0.06fF
C60 w_1856_392# OUT6 0.06fF
C61 VDD OUT8 0.21fF
C62 OUT7 Gnd 0.14fF
C63 In6 a_1777_355# 0.19fF
C64 VDD OUT7 0.21fF
C65 OUT6 Gnd 0.14fF
C66 a_1561_407# a_1574_355# 0.21fF
C67 In3 a_1156_407# 0.10fF
C68 VDD OUT6 0.21fF
C69 OUT5 Gnd 0.14fF
C70 In1 a_766_407# 0.10fF
C71 w_1450_392# a_1358_407# 0.06fF
C72 VDD OUT5 0.21fF
C73 OUT4 Gnd 0.14fF
C74 In2 a_964_407# 0.10fF
C75 VDD OUT4 0.21fF
C76 w_1248_392# OUT3 0.06fF
C77 OUT3 Gnd 0.14fF
C78 In3 a_1169_355# 0.19fF
C79 VDD OUT3 0.21fF
C80 OUT2 Gnd 0.14fF
C81 a_964_407# a_977_355# 0.21fF
C82 w_858_392# a_766_407# 0.06fF
C83 In1 a_779_355# 0.19fF
C84 Gnd a_1981_355# 0.21fF
C85 VDD OUT2 0.21fF
C86 w_858_392# OUT1 0.06fF
C87 VDD EN 21.53fF
C88 EN a_2171_407# 0.47fF
C89 w_2263_392# OUT8 0.06fF
C90 Gnd a_1371_355# 0.21fF
C91 In8 a_2184_355# 0.19fF
C92 VDD w_1856_392# 0.06fF
C93 EN a_1968_407# 0.47fF
C94 a_1968_407# a_1981_355# 0.21fF
C95 VDD w_1248_392# 0.06fF
C96 EN a_1764_407# 0.47fF
C97 a_2184_355# Gnd 0.20fF
C98 a_1981_355# Gnd 0.20fF
C99 a_1777_355# Gnd 0.20fF
C100 a_1574_355# Gnd 0.20fF
C101 a_1371_355# Gnd 0.20fF
C102 a_1169_355# Gnd 0.20fF
C103 a_977_355# Gnd 0.20fF
C104 Gnd Gnd 0.32fF
C105 a_779_355# Gnd 0.20fF
C106 OUT8 Gnd 0.13fF
C107 a_2171_407# Gnd 0.78fF
C108 In8 Gnd 0.49fF
C109 OUT7 Gnd 0.13fF
C110 a_1968_407# Gnd 0.78fF
C111 In7 Gnd 0.49fF
C112 OUT6 Gnd 0.13fF
C113 a_1764_407# Gnd 0.78fF
C114 In6 Gnd 0.49fF
C115 OUT5 Gnd 0.13fF
C116 a_1561_407# Gnd 0.78fF
C117 In5 Gnd 0.49fF
C118 OUT4 Gnd 0.13fF
C119 a_1358_407# Gnd 0.78fF
C120 In4 Gnd 0.49fF
C121 OUT3 Gnd 0.13fF
C122 a_1156_407# Gnd 0.78fF
C123 In3 Gnd 0.49fF
C124 OUT2 Gnd 0.13fF
C125 a_964_407# Gnd 0.78fF
C126 In2 Gnd 0.49fF
C127 OUT1 Gnd 0.13fF
C128 a_766_407# Gnd 0.78fF
C129 In1 Gnd 0.99fF
C130 EN Gnd 0.62fF
C131 w_2263_392# Gnd 1.16fF
C132 w_2060_392# Gnd 1.16fF
C133 w_1856_392# Gnd 1.16fF
C134 w_1653_392# Gnd 1.16fF
C135 w_1450_392# Gnd 1.16fF
C136 w_1248_392# Gnd 1.16fF
C137 w_1056_392# Gnd 1.16fF
C138 w_858_392# Gnd 1.16fF
C139 VDD Gnd 23.05fF

.tran 1n 10n
.control
run
set color0 = white
set color1 = black
plot v(OUT1) v(OUT2)+2 v(OUT3)+4 v(OUT4)+6 v(OUT5)+8 v(OUT6)+10 v(OUT7)+12 v(OUT8)+14 v(EN)+16
.endc
.end