magic
tech scmos
timestamp 1701501258
<< nwell >>
rect 278 174 314 206
rect 334 174 370 206
rect 390 174 426 206
rect 446 174 482 206
rect 501 174 537 206
<< ntransistor >>
rect 321 128 325 148
rect 321 88 325 108
rect 321 48 325 68
rect 321 9 325 29
rect 321 -30 325 -10
<< ptransistor >>
rect 295 180 297 200
rect 351 180 353 200
rect 407 180 409 200
rect 463 180 465 200
rect 518 180 520 200
<< ndiffusion >>
rect 320 128 321 148
rect 325 128 326 148
rect 320 88 321 108
rect 325 88 326 108
rect 320 48 321 68
rect 325 48 326 68
rect 320 9 321 29
rect 325 9 326 29
rect 320 -30 321 -10
rect 325 -30 326 -10
<< pdiffusion >>
rect 294 180 295 200
rect 297 180 298 200
rect 350 180 351 200
rect 353 180 354 200
rect 406 180 407 200
rect 409 180 410 200
rect 462 180 463 200
rect 465 180 466 200
rect 517 180 518 200
rect 520 180 521 200
<< ndcontact >>
rect 310 128 320 148
rect 326 128 336 148
rect 310 88 320 108
rect 326 88 336 108
rect 310 48 320 68
rect 326 48 336 68
rect 310 9 320 29
rect 326 9 336 29
rect 310 -30 320 -10
rect 326 -30 336 -10
<< pdcontact >>
rect 284 180 294 200
rect 298 180 308 200
rect 340 180 350 200
rect 354 180 364 200
rect 396 180 406 200
rect 410 180 420 200
rect 452 180 462 200
rect 466 180 476 200
rect 507 180 517 200
rect 521 180 531 200
<< psubstratepcontact >>
rect 278 -39 282 -35
rect 533 -39 537 -35
<< nsubstratencontact >>
rect 278 206 282 210
rect 533 206 537 210
<< polysilicon >>
rect 295 200 297 203
rect 351 200 353 203
rect 407 200 409 203
rect 463 200 465 203
rect 518 200 520 203
rect 295 171 297 180
rect 351 171 353 180
rect 407 171 409 180
rect 463 171 465 180
rect 518 171 520 180
rect 282 167 297 171
rect 338 167 353 171
rect 394 167 409 171
rect 450 167 465 171
rect 505 167 520 171
rect 310 151 325 155
rect 321 148 325 151
rect 321 125 325 128
rect 349 115 353 167
rect 310 111 353 115
rect 321 108 325 111
rect 321 85 325 88
rect 405 75 409 167
rect 310 71 409 75
rect 321 68 325 71
rect 321 45 325 48
rect 461 36 465 167
rect 310 32 465 36
rect 321 29 325 32
rect 321 6 325 9
rect 516 -3 520 167
rect 310 -7 520 -3
rect 321 -10 325 -7
rect 321 -33 325 -30
<< polycontact >>
rect 278 167 282 171
rect 306 151 310 155
rect 306 111 310 115
rect 306 71 310 75
rect 306 32 310 36
rect 306 -7 310 -3
<< metal1 >>
rect 282 206 533 210
rect 284 200 294 206
rect 340 200 350 206
rect 396 200 406 206
rect 452 200 462 206
rect 507 200 517 206
rect 263 167 278 171
rect 263 155 267 167
rect 298 162 308 180
rect 354 162 364 180
rect 410 162 420 180
rect 466 162 476 180
rect 521 162 531 180
rect 278 158 537 162
rect 263 151 306 155
rect 326 148 336 158
rect 310 122 320 128
rect 310 118 336 122
rect 291 111 306 115
rect 326 108 336 118
rect 310 82 320 88
rect 310 78 336 82
rect 291 71 306 75
rect 326 68 336 78
rect 310 43 320 48
rect 310 39 336 43
rect 291 32 306 36
rect 326 29 336 39
rect 310 4 320 9
rect 310 0 336 4
rect 291 -7 306 -3
rect 326 -10 336 0
rect 310 -35 320 -30
rect 282 -39 533 -35
<< labels >>
rlabel metal1 263 167 282 171 1 A
rlabel metal1 291 111 310 115 1 B
rlabel metal1 291 71 310 75 1 C
rlabel metal1 291 32 310 36 1 D
rlabel metal1 278 -39 537 -35 1 Gnd
rlabel metal1 278 158 537 162 1 OUT
rlabel metal1 278 206 537 210 5 VDD
rlabel metal1 291 -7 310 -3 1 E
<< end >>
