ARITHMATIC_LOGIC_UNIT 4 Bit

* Technology File
.include TSMC_180nm.txt

* Gates Required
.include AND2.sub
.include AND3.sub
.include AND4.sub
.include NAND2.sub
.include NAND3.sub
.include NAND4.sub
.include NAND5.sub
.include NOR2.sub
.include NOT.sub
.include OR2.sub
.include XNOR2.sub
.include XOR2.sub

* Component Subcircuits
.include decoder.sub
.include Enable.sub
.include FA.sub
.include adder_subtractor.sub
.include comparator.sub
.include and_4bit.sub

.param SUPPLY = 1.8
.param LAMBDA = 0.18u

* Width and Length of NMOS
.param wn1 = {10*LAMBDA}
.param ln1 = {2*LAMBDA}
.param wn2 = {10*LAMBDA}
.param ln2 = {2*LAMBDA}
.param wn3 = {10*LAMBDA}
.param ln3 = {2*LAMBDA}
.param wn4 = {10*LAMBDA}
.param ln4 = {2*LAMBDA}
.param wn5 = {10*LAMBDA}
.param ln5 = {2*LAMBDA}

* Width and Length of NMOS
.param wp1 = wn1
.param lp1 = {LAMBDA}
.param wp2 = wn2
.param lp2 = {LAMBDA}
.param wp3 = wn3
.param lp3 = {LAMBDA}
.param wp4 = wn4
.param lp4 = {LAMBDA}
.param wp5 = wn5
.param lp5 = {LAMBDA}

.global GND

Vdd V GND 'SUPPLY'

VS0 S0 Gnd DC 'SUPPLY'
VS1 S1 Gnd DC 0

VA3 A3 Gnd DC 1
VA2 A2 Gnd DC 1
VA1 A1 Gnd DC 1
VA0 A0 Gnd DC 1

VB3 B3 Gnd PULSE('SUPPLY' 0 0ns 100ps 100ps 10ns 20ns)
VB2 B2 Gnd PULSE('SUPPLY' 0 0ns 100ps 100ps 10ns 20ns)
VB1 B1 Gnd PULSE('SUPPLY' 0 0ns 100ps 100ps 10ns 20ns)
VB0 B0 Gnd PULSE('SUPPLY' 0 0ns 100ps 100ps 10ns 20ns)

* Decode based on select lines
X_DEC S1 S0 D0 D1 D2 D3 V GND decoder
*Adder/Subtractor
X_R2 D0 D1 DAS V GND OR2
X_EN1 A3 A2 A1 A0 B3 B2 B1 B0 DAS ASA3 ASA2 ASA1 ASA0 ASB3 ASB2 ASB1 ASB0 V GND Enable
X_AS ASA3 ASA2 ASA1 ASA0 ASB3 ASB2 ASB1 ASB0 D1 C OUT_AS3 OUT_AS2 OUT_AS1 OUT_AS0 V GND adder_subtractor
*Comparator
X_EN2 A3 A2 A1 A0 B3 B2 B1 B0 D2 COA3 COA2 COA1 COA0 COB3 COB2 COB1 COB0 V GND Enable
X_COMP COA3 COA2 COA1 COA0 COB3 COB2 COB1 COB0 E1 G L V GND comparator
X_And2 E1 D2 E V GND AND2
* 4 Bit And
X_EN3 A3 A2 A1 A0 B3 B2 B1 B0 D3 ANA3 ANA2 ANA1 ANA0 ANB3 ANB2 ANB1 ANB0 V GND Enable
X_AN ANA3 ANA2 ANA1 ANA0 ANB3 ANB2 ANB1 ANB0 OUT_AND3 OUT_AND2 OUT_AND1 OUT_AND0 V GND and_4bit

.tran 1n 80n


.measure tran trise 
+ TRIG v(B3) VAL = 'SUPPLY/2' RISE =1
+ TARG v(E) VAL = 'SUPPLY/2' RISE =1 

.measure tran tfall 
+ TRIG v(B3) VAL = 'SUPPLY/2' FALL =1 
+ TARG v(E) VAL = 'SUPPLY/2' FALL=1

.measure tran tpd param = '(trise + tfall)/2' goal = 0


.control 

    run
    quit

.endc
.end
