module and_4bit_tb;
    reg A3,A2,A1,A0,B3,B2,B0,B1;
    wire out3,out2,out1,out0;

    and_4bit and_4bit_tb(A3,A2,A1,A0,B3,B2,B1,B0,out3,out2,out1,out0);
    initial
    begin
        $dumpfile("and_4bit_out.vcd");
        $dumpvars(0,and_4bit_tb);
        $monitor("T=%4t:A3 = %b,A2 = %b,A1 = %b,A0 = %b,B3 = %b,B2 = %b,B1 = %b,B0 = %b, out3 = %b, out2 = %b, out1 = %b, out0 = %b",$time,A3,A2,A1,A0,B3,B2,B1,B0,out3,out2,out1,out0);
        #5 A3=0;A2=0;A1=0;A0=0;B3=0;B2=0;B1=0;B0=0;
        #5 A3=0;A2=0;A1=0;A0=0;B3=0;B2=0;B1=0;B0=1;
        #5 A3=0;A2=0;A1=0;A0=0;B3=0;B2=0;B1=1;B0=0;
        #5 A3=0;A2=0;A1=0;A0=0;B3=0;B2=0;B1=1;B0=1;
        #5 A3=0;A2=0;A1=0;A0=0;B3=0;B2=1;B1=0;B0=0;
        #5 A3=0;A2=0;A1=0;A0=0;B3=0;B2=1;B1=0;B0=1;
        #5 A3=0;A2=0;A1=0;A0=0;B3=0;B2=1;B1=1;B0=0;
        #5 A3=0;A2=0;A1=0;A0=0;B3=0;B2=1;B1=1;B0=1;
        #5 A3=0;A2=0;A1=0;A0=0;B3=1;B2=0;B1=0;B0=0;
        #5 A3=0;A2=0;A1=0;A0=0;B3=1;B2=0;B1=0;B0=1;
        #5 A3=0;A2=0;A1=0;A0=0;B3=1;B2=0;B1=1;B0=0;
        #5 A3=0;A2=0;A1=0;A0=0;B3=1;B2=0;B1=1;B0=1;
        #5 A3=0;A2=0;A1=0;A0=0;B3=1;B2=1;B1=0;B0=0;
        #5 A3=0;A2=0;A1=0;A0=0;B3=1;B2=1;B1=0;B0=1;
        #5 A3=0;A2=0;A1=0;A0=0;B3=1;B2=1;B1=1;B0=0;
        #5 A3=0;A2=0;A1=0;A0=0;B3=1;B2=1;B1=1;B0=1;
        #5 A3=0;A2=0;A1=0;A0=1;B3=0;B2=0;B1=0;B0=0;
        #5 A3=0;A2=0;A1=0;A0=1;B3=0;B2=0;B1=0;B0=1;
        #5 A3=0;A2=0;A1=0;A0=1;B3=0;B2=0;B1=1;B0=0;
        #5 A3=0;A2=0;A1=0;A0=1;B3=0;B2=0;B1=1;B0=1;
        #5 A3=0;A2=0;A1=0;A0=1;B3=0;B2=1;B1=0;B0=0;
        #5 A3=0;A2=0;A1=0;A0=1;B3=0;B2=1;B1=0;B0=1;
        #5 A3=0;A2=0;A1=0;A0=1;B3=0;B2=1;B1=1;B0=0;
        #5 A3=0;A2=0;A1=0;A0=1;B3=0;B2=1;B1=1;B0=1;
        #5 A3=0;A2=0;A1=0;A0=1;B3=1;B2=0;B1=0;B0=0;
        #5 A3=0;A2=0;A1=0;A0=1;B3=1;B2=0;B1=0;B0=1;
        #5 A3=0;A2=0;A1=0;A0=1;B3=1;B2=0;B1=1;B0=0;
        #5 A3=0;A2=0;A1=0;A0=1;B3=1;B2=0;B1=1;B0=1;
        #5 A3=0;A2=0;A1=0;A0=1;B3=1;B2=1;B1=0;B0=0;
        #5 A3=0;A2=0;A1=0;A0=1;B3=1;B2=1;B1=0;B0=1;
        #5 A3=0;A2=0;A1=0;A0=1;B3=1;B2=1;B1=1;B0=0;
        #5 A3=0;A2=0;A1=0;A0=1;B3=1;B2=1;B1=1;B0=1;
        #5 A3=0;A2=0;A1=1;A0=0;B3=0;B2=0;B1=0;B0=0;
        #5 A3=0;A2=0;A1=1;A0=0;B3=0;B2=0;B1=0;B0=1;
        #5 A3=0;A2=0;A1=1;A0=0;B3=0;B2=0;B1=1;B0=0;
        #5 A3=0;A2=0;A1=1;A0=0;B3=0;B2=0;B1=1;B0=1;
        #5 A3=0;A2=0;A1=1;A0=0;B3=0;B2=1;B1=0;B0=0;
        #5 A3=0;A2=0;A1=1;A0=0;B3=0;B2=1;B1=0;B0=1;
        #5 A3=0;A2=0;A1=1;A0=0;B3=0;B2=1;B1=1;B0=0;
        #5 A3=0;A2=0;A1=1;A0=0;B3=0;B2=1;B1=1;B0=1;
        #5 A3=0;A2=0;A1=1;A0=0;B3=1;B2=0;B1=0;B0=0;
        #5 A3=0;A2=0;A1=1;A0=0;B3=1;B2=0;B1=0;B0=1;
        #5 A3=0;A2=0;A1=1;A0=0;B3=1;B2=0;B1=1;B0=0;
        #5 A3=0;A2=0;A1=1;A0=0;B3=1;B2=0;B1=1;B0=1;
        #5 A3=0;A2=0;A1=1;A0=0;B3=1;B2=1;B1=0;B0=0;
        #5 A3=0;A2=0;A1=1;A0=0;B3=1;B2=1;B1=0;B0=1;
        #5 A3=0;A2=0;A1=1;A0=0;B3=1;B2=1;B1=1;B0=0;
        #5 A3=0;A2=0;A1=1;A0=0;B3=1;B2=1;B1=1;B0=1;
        #5 A3=0;A2=0;A1=1;A0=1;B3=0;B2=0;B1=0;B0=0;
        #5 A3=0;A2=0;A1=1;A0=1;B3=0;B2=0;B1=0;B0=1;
        #5 A3=0;A2=0;A1=1;A0=1;B3=0;B2=0;B1=1;B0=0;
        #5 A3=0;A2=0;A1=1;A0=1;B3=0;B2=0;B1=1;B0=1;
        #5 A3=0;A2=0;A1=1;A0=1;B3=0;B2=1;B1=0;B0=0;
        #5 A3=0;A2=0;A1=1;A0=1;B3=0;B2=1;B1=0;B0=1;
        #5 A3=0;A2=0;A1=1;A0=1;B3=0;B2=1;B1=1;B0=0;
        #5 A3=0;A2=0;A1=1;A0=1;B3=0;B2=1;B1=1;B0=1;
        #5 A3=0;A2=0;A1=1;A0=1;B3=1;B2=0;B1=0;B0=0;
        #5 A3=0;A2=0;A1=1;A0=1;B3=1;B2=0;B1=0;B0=1;
        #5 A3=0;A2=0;A1=1;A0=1;B3=1;B2=0;B1=1;B0=0;
        #5 A3=0;A2=0;A1=1;A0=1;B3=1;B2=0;B1=1;B0=1;
        #5 A3=0;A2=0;A1=1;A0=1;B3=1;B2=1;B1=0;B0=0;
        #5 A3=0;A2=0;A1=1;A0=1;B3=1;B2=1;B1=0;B0=1;
        #5 A3=0;A2=0;A1=1;A0=1;B3=1;B2=1;B1=1;B0=0;
        #5 A3=0;A2=0;A1=1;A0=1;B3=1;B2=1;B1=1;B0=1;
        #5 A3=0;A2=1;A1=0;A0=0;B3=0;B2=0;B1=0;B0=0;
        #5 A3=0;A2=1;A1=0;A0=0;B3=0;B2=0;B1=0;B0=1;
        #5 A3=0;A2=1;A1=0;A0=0;B3=0;B2=0;B1=1;B0=0;
        #5 A3=0;A2=1;A1=0;A0=0;B3=0;B2=0;B1=1;B0=1;
        #5 A3=0;A2=1;A1=0;A0=0;B3=0;B2=1;B1=0;B0=0;
        #5 A3=0;A2=1;A1=0;A0=0;B3=0;B2=1;B1=0;B0=1;
        #5 A3=0;A2=1;A1=0;A0=0;B3=0;B2=1;B1=1;B0=0;
        #5 A3=0;A2=1;A1=0;A0=0;B3=0;B2=1;B1=1;B0=1;
        #5 A3=0;A2=1;A1=0;A0=0;B3=1;B2=0;B1=0;B0=0;
        #5 A3=0;A2=1;A1=0;A0=0;B3=1;B2=0;B1=0;B0=1;
        #5 A3=0;A2=1;A1=0;A0=0;B3=1;B2=0;B1=1;B0=0;
        #5 A3=0;A2=1;A1=0;A0=0;B3=1;B2=0;B1=1;B0=1;
        #5 A3=0;A2=1;A1=0;A0=0;B3=1;B2=1;B1=0;B0=0;
        #5 A3=0;A2=1;A1=0;A0=0;B3=1;B2=1;B1=0;B0=1;
        #5 A3=0;A2=1;A1=0;A0=0;B3=1;B2=1;B1=1;B0=0;
        #5 A3=0;A2=1;A1=0;A0=0;B3=1;B2=1;B1=1;B0=1;
        #5 A3=0;A2=1;A1=0;A0=1;B3=0;B2=0;B1=0;B0=0;
        #5 A3=0;A2=1;A1=0;A0=1;B3=0;B2=0;B1=0;B0=1;
        #5 A3=0;A2=1;A1=0;A0=1;B3=0;B2=0;B1=1;B0=0;
        #5 A3=0;A2=1;A1=0;A0=1;B3=0;B2=0;B1=1;B0=1;
        #5 A3=0;A2=1;A1=0;A0=1;B3=0;B2=1;B1=0;B0=0;
        #5 A3=0;A2=1;A1=0;A0=1;B3=0;B2=1;B1=0;B0=1;
        #5 A3=0;A2=1;A1=0;A0=1;B3=0;B2=1;B1=1;B0=0;
        #5 A3=0;A2=1;A1=0;A0=1;B3=0;B2=1;B1=1;B0=1;
        #5 A3=0;A2=1;A1=0;A0=1;B3=1;B2=0;B1=0;B0=0;
        #5 A3=0;A2=1;A1=0;A0=1;B3=1;B2=0;B1=0;B0=1;
        #5 A3=0;A2=1;A1=0;A0=1;B3=1;B2=0;B1=1;B0=0;
        #5 A3=0;A2=1;A1=0;A0=1;B3=1;B2=0;B1=1;B0=1;
        #5 A3=0;A2=1;A1=0;A0=1;B3=1;B2=1;B1=0;B0=0;
        #5 A3=0;A2=1;A1=0;A0=1;B3=1;B2=1;B1=0;B0=1;
        #5 A3=0;A2=1;A1=0;A0=1;B3=1;B2=1;B1=1;B0=0;
        #5 A3=0;A2=1;A1=0;A0=1;B3=1;B2=1;B1=1;B0=1;
        #5 A3=0;A2=1;A1=1;A0=0;B3=0;B2=0;B1=0;B0=0;
        #5 A3=0;A2=1;A1=1;A0=0;B3=0;B2=0;B1=0;B0=1;
        #5 A3=0;A2=1;A1=1;A0=0;B3=0;B2=0;B1=1;B0=0;
        #5 A3=0;A2=1;A1=1;A0=0;B3=0;B2=0;B1=1;B0=1;
        #5 A3=0;A2=1;A1=1;A0=0;B3=0;B2=1;B1=0;B0=0;
        #5 A3=0;A2=1;A1=1;A0=0;B3=0;B2=1;B1=0;B0=1;
        #5 A3=0;A2=1;A1=1;A0=0;B3=0;B2=1;B1=1;B0=0;
        #5 A3=0;A2=1;A1=1;A0=0;B3=0;B2=1;B1=1;B0=1;
        #5 A3=0;A2=1;A1=1;A0=0;B3=1;B2=0;B1=0;B0=0;
        #5 A3=0;A2=1;A1=1;A0=0;B3=1;B2=0;B1=0;B0=1;
        #5 A3=0;A2=1;A1=1;A0=0;B3=1;B2=0;B1=1;B0=0;
        #5 A3=0;A2=1;A1=1;A0=0;B3=1;B2=0;B1=1;B0=1;
        #5 A3=0;A2=1;A1=1;A0=0;B3=1;B2=1;B1=0;B0=0;
        #5 A3=0;A2=1;A1=1;A0=0;B3=1;B2=1;B1=0;B0=1;
        #5 A3=0;A2=1;A1=1;A0=0;B3=1;B2=1;B1=1;B0=0;
        #5 A3=0;A2=1;A1=1;A0=0;B3=1;B2=1;B1=1;B0=1;
        #5 A3=0;A2=1;A1=1;A0=1;B3=0;B2=0;B1=0;B0=0;
        #5 A3=0;A2=1;A1=1;A0=1;B3=0;B2=0;B1=0;B0=1;
        #5 A3=0;A2=1;A1=1;A0=1;B3=0;B2=0;B1=1;B0=0;
        #5 A3=0;A2=1;A1=1;A0=1;B3=0;B2=0;B1=1;B0=1;
        #5 A3=0;A2=1;A1=1;A0=1;B3=0;B2=1;B1=0;B0=0;
        #5 A3=0;A2=1;A1=1;A0=1;B3=0;B2=1;B1=0;B0=1;
        #5 A3=0;A2=1;A1=1;A0=1;B3=0;B2=1;B1=1;B0=0;
        #5 A3=0;A2=1;A1=1;A0=1;B3=0;B2=1;B1=1;B0=1;
        #5 A3=0;A2=1;A1=1;A0=1;B3=1;B2=0;B1=0;B0=0;
        #5 A3=0;A2=1;A1=1;A0=1;B3=1;B2=0;B1=0;B0=1;
        #5 A3=0;A2=1;A1=1;A0=1;B3=1;B2=0;B1=1;B0=0;
        #5 A3=0;A2=1;A1=1;A0=1;B3=1;B2=0;B1=1;B0=1;
        #5 A3=0;A2=1;A1=1;A0=1;B3=1;B2=1;B1=0;B0=0;
        #5 A3=0;A2=1;A1=1;A0=1;B3=1;B2=1;B1=0;B0=1;
        #5 A3=0;A2=1;A1=1;A0=1;B3=1;B2=1;B1=1;B0=0;
        #5 A3=0;A2=1;A1=1;A0=1;B3=1;B2=1;B1=1;B0=1;
        #5 A3=1;A2=0;A1=0;A0=0;B3=0;B2=0;B1=0;B0=0;
        #5 A3=1;A2=0;A1=0;A0=0;B3=0;B2=0;B1=0;B0=1;
        #5 A3=1;A2=0;A1=0;A0=0;B3=0;B2=0;B1=1;B0=0;
        #5 A3=1;A2=0;A1=0;A0=0;B3=0;B2=0;B1=1;B0=1;
        #5 A3=1;A2=0;A1=0;A0=0;B3=0;B2=1;B1=0;B0=0;
        #5 A3=1;A2=0;A1=0;A0=0;B3=0;B2=1;B1=0;B0=1;
        #5 A3=1;A2=0;A1=0;A0=0;B3=0;B2=1;B1=1;B0=0;
        #5 A3=1;A2=0;A1=0;A0=0;B3=0;B2=1;B1=1;B0=1;
        #5 A3=1;A2=0;A1=0;A0=0;B3=1;B2=0;B1=0;B0=0;
        #5 A3=1;A2=0;A1=0;A0=0;B3=1;B2=0;B1=0;B0=1;
        #5 A3=1;A2=0;A1=0;A0=0;B3=1;B2=0;B1=1;B0=0;
        #5 A3=1;A2=0;A1=0;A0=0;B3=1;B2=0;B1=1;B0=1;
        #5 A3=1;A2=0;A1=0;A0=0;B3=1;B2=1;B1=0;B0=0;
        #5 A3=1;A2=0;A1=0;A0=0;B3=1;B2=1;B1=0;B0=1;
        #5 A3=1;A2=0;A1=0;A0=0;B3=1;B2=1;B1=1;B0=0;
        #5 A3=1;A2=0;A1=0;A0=0;B3=1;B2=1;B1=1;B0=1;
        #5 A3=1;A2=0;A1=0;A0=1;B3=0;B2=0;B1=0;B0=0;
        #5 A3=1;A2=0;A1=0;A0=1;B3=0;B2=0;B1=0;B0=1;
        #5 A3=1;A2=0;A1=0;A0=1;B3=0;B2=0;B1=1;B0=0;
        #5 A3=1;A2=0;A1=0;A0=1;B3=0;B2=0;B1=1;B0=1;
        #5 A3=1;A2=0;A1=0;A0=1;B3=0;B2=1;B1=0;B0=0;
        #5 A3=1;A2=0;A1=0;A0=1;B3=0;B2=1;B1=0;B0=1;
        #5 A3=1;A2=0;A1=0;A0=1;B3=0;B2=1;B1=1;B0=0;
        #5 A3=1;A2=0;A1=0;A0=1;B3=0;B2=1;B1=1;B0=1;
        #5 A3=1;A2=0;A1=0;A0=1;B3=1;B2=0;B1=0;B0=0;
        #5 A3=1;A2=0;A1=0;A0=1;B3=1;B2=0;B1=0;B0=1;
        #5 A3=1;A2=0;A1=0;A0=1;B3=1;B2=0;B1=1;B0=0;
        #5 A3=1;A2=0;A1=0;A0=1;B3=1;B2=0;B1=1;B0=1;
        #5 A3=1;A2=0;A1=0;A0=1;B3=1;B2=1;B1=0;B0=0;
        #5 A3=1;A2=0;A1=0;A0=1;B3=1;B2=1;B1=0;B0=1;
        #5 A3=1;A2=0;A1=0;A0=1;B3=1;B2=1;B1=1;B0=0;
        #5 A3=1;A2=0;A1=0;A0=1;B3=1;B2=1;B1=1;B0=1;
        #5 A3=1;A2=0;A1=1;A0=0;B3=0;B2=0;B1=0;B0=0;
        #5 A3=1;A2=0;A1=1;A0=0;B3=0;B2=0;B1=0;B0=1;
        #5 A3=1;A2=0;A1=1;A0=0;B3=0;B2=0;B1=1;B0=0;
        #5 A3=1;A2=0;A1=1;A0=0;B3=0;B2=0;B1=1;B0=1;
        #5 A3=1;A2=0;A1=1;A0=0;B3=0;B2=1;B1=0;B0=0;
        #5 A3=1;A2=0;A1=1;A0=0;B3=0;B2=1;B1=0;B0=1;
        #5 A3=1;A2=0;A1=1;A0=0;B3=0;B2=1;B1=1;B0=0;
        #5 A3=1;A2=0;A1=1;A0=0;B3=0;B2=1;B1=1;B0=1;
        #5 A3=1;A2=0;A1=1;A0=0;B3=1;B2=0;B1=0;B0=0;
        #5 A3=1;A2=0;A1=1;A0=0;B3=1;B2=0;B1=0;B0=1;
        #5 A3=1;A2=0;A1=1;A0=0;B3=1;B2=0;B1=1;B0=0;
        #5 A3=1;A2=0;A1=1;A0=0;B3=1;B2=0;B1=1;B0=1;
        #5 A3=1;A2=0;A1=1;A0=0;B3=1;B2=1;B1=0;B0=0;
        #5 A3=1;A2=0;A1=1;A0=0;B3=1;B2=1;B1=0;B0=1;
        #5 A3=1;A2=0;A1=1;A0=0;B3=1;B2=1;B1=1;B0=0;
        #5 A3=1;A2=0;A1=1;A0=0;B3=1;B2=1;B1=1;B0=1;
        #5 A3=1;A2=0;A1=1;A0=1;B3=0;B2=0;B1=0;B0=0;
        #5 A3=1;A2=0;A1=1;A0=1;B3=0;B2=0;B1=0;B0=1;
        #5 A3=1;A2=0;A1=1;A0=1;B3=0;B2=0;B1=1;B0=0;
        #5 A3=1;A2=0;A1=1;A0=1;B3=0;B2=0;B1=1;B0=1;
        #5 A3=1;A2=0;A1=1;A0=1;B3=0;B2=1;B1=0;B0=0;
        #5 A3=1;A2=0;A1=1;A0=1;B3=0;B2=1;B1=0;B0=1;
        #5 A3=1;A2=0;A1=1;A0=1;B3=0;B2=1;B1=1;B0=0;
        #5 A3=1;A2=0;A1=1;A0=1;B3=0;B2=1;B1=1;B0=1;
        #5 A3=1;A2=0;A1=1;A0=1;B3=1;B2=0;B1=0;B0=0;
        #5 A3=1;A2=0;A1=1;A0=1;B3=1;B2=0;B1=0;B0=1;
        #5 A3=1;A2=0;A1=1;A0=1;B3=1;B2=0;B1=1;B0=0;
        #5 A3=1;A2=0;A1=1;A0=1;B3=1;B2=0;B1=1;B0=1;
        #5 A3=1;A2=0;A1=1;A0=1;B3=1;B2=1;B1=0;B0=0;
        #5 A3=1;A2=0;A1=1;A0=1;B3=1;B2=1;B1=0;B0=1;
        #5 A3=1;A2=0;A1=1;A0=1;B3=1;B2=1;B1=1;B0=0;
        #5 A3=1;A2=0;A1=1;A0=1;B3=1;B2=1;B1=1;B0=1;
        #5 A3=1;A2=1;A1=0;A0=0;B3=0;B2=0;B1=0;B0=0;
        #5 A3=1;A2=1;A1=0;A0=0;B3=0;B2=0;B1=0;B0=1;
        #5 A3=1;A2=1;A1=0;A0=0;B3=0;B2=0;B1=1;B0=0;
        #5 A3=1;A2=1;A1=0;A0=0;B3=0;B2=0;B1=1;B0=1;
        #5 A3=1;A2=1;A1=0;A0=0;B3=0;B2=1;B1=0;B0=0;
        #5 A3=1;A2=1;A1=0;A0=0;B3=0;B2=1;B1=0;B0=1;
        #5 A3=1;A2=1;A1=0;A0=0;B3=0;B2=1;B1=1;B0=0;
        #5 A3=1;A2=1;A1=0;A0=0;B3=0;B2=1;B1=1;B0=1;
        #5 A3=1;A2=1;A1=0;A0=0;B3=1;B2=0;B1=0;B0=0;
        #5 A3=1;A2=1;A1=0;A0=0;B3=1;B2=0;B1=0;B0=1;
        #5 A3=1;A2=1;A1=0;A0=0;B3=1;B2=0;B1=1;B0=0;
        #5 A3=1;A2=1;A1=0;A0=0;B3=1;B2=0;B1=1;B0=1;
        #5 A3=1;A2=1;A1=0;A0=0;B3=1;B2=1;B1=0;B0=0;
        #5 A3=1;A2=1;A1=0;A0=0;B3=1;B2=1;B1=0;B0=1;
        #5 A3=1;A2=1;A1=0;A0=0;B3=1;B2=1;B1=1;B0=0;
        #5 A3=1;A2=1;A1=0;A0=0;B3=1;B2=1;B1=1;B0=1;
        #5 A3=1;A2=1;A1=0;A0=1;B3=0;B2=0;B1=0;B0=0;
        #5 A3=1;A2=1;A1=0;A0=1;B3=0;B2=0;B1=0;B0=1;
        #5 A3=1;A2=1;A1=0;A0=1;B3=0;B2=0;B1=1;B0=0;
        #5 A3=1;A2=1;A1=0;A0=1;B3=0;B2=0;B1=1;B0=1;
        #5 A3=1;A2=1;A1=0;A0=1;B3=0;B2=1;B1=0;B0=0;
        #5 A3=1;A2=1;A1=0;A0=1;B3=0;B2=1;B1=0;B0=1;
        #5 A3=1;A2=1;A1=0;A0=1;B3=0;B2=1;B1=1;B0=0;
        #5 A3=1;A2=1;A1=0;A0=1;B3=0;B2=1;B1=1;B0=1;
        #5 A3=1;A2=1;A1=0;A0=1;B3=1;B2=0;B1=0;B0=0;
        #5 A3=1;A2=1;A1=0;A0=1;B3=1;B2=0;B1=0;B0=1;
        #5 A3=1;A2=1;A1=0;A0=1;B3=1;B2=0;B1=1;B0=0;
        #5 A3=1;A2=1;A1=0;A0=1;B3=1;B2=0;B1=1;B0=1;
        #5 A3=1;A2=1;A1=0;A0=1;B3=1;B2=1;B1=0;B0=0;
        #5 A3=1;A2=1;A1=0;A0=1;B3=1;B2=1;B1=0;B0=1;
        #5 A3=1;A2=1;A1=0;A0=1;B3=1;B2=1;B1=1;B0=0;
        #5 A3=1;A2=1;A1=0;A0=1;B3=1;B2=1;B1=1;B0=1;
        #5 A3=1;A2=1;A1=1;A0=0;B3=0;B2=0;B1=0;B0=0;
        #5 A3=1;A2=1;A1=1;A0=0;B3=0;B2=0;B1=0;B0=1;
        #5 A3=1;A2=1;A1=1;A0=0;B3=0;B2=0;B1=1;B0=0;
        #5 A3=1;A2=1;A1=1;A0=0;B3=0;B2=0;B1=1;B0=1;
        #5 A3=1;A2=1;A1=1;A0=0;B3=0;B2=1;B1=0;B0=0;
        #5 A3=1;A2=1;A1=1;A0=0;B3=0;B2=1;B1=0;B0=1;
        #5 A3=1;A2=1;A1=1;A0=0;B3=0;B2=1;B1=1;B0=0;
        #5 A3=1;A2=1;A1=1;A0=0;B3=0;B2=1;B1=1;B0=1;
        #5 A3=1;A2=1;A1=1;A0=0;B3=1;B2=0;B1=0;B0=0;
        #5 A3=1;A2=1;A1=1;A0=0;B3=1;B2=0;B1=0;B0=1;
        #5 A3=1;A2=1;A1=1;A0=0;B3=1;B2=0;B1=1;B0=0;
        #5 A3=1;A2=1;A1=1;A0=0;B3=1;B2=0;B1=1;B0=1;
        #5 A3=1;A2=1;A1=1;A0=0;B3=1;B2=1;B1=0;B0=0;
        #5 A3=1;A2=1;A1=1;A0=0;B3=1;B2=1;B1=0;B0=1;
        #5 A3=1;A2=1;A1=1;A0=0;B3=1;B2=1;B1=1;B0=0;
        #5 A3=1;A2=1;A1=1;A0=0;B3=1;B2=1;B1=1;B0=1;
        #5 A3=1;A2=1;A1=1;A0=1;B3=0;B2=0;B1=0;B0=0;
        #5 A3=1;A2=1;A1=1;A0=1;B3=0;B2=0;B1=0;B0=1;
        #5 A3=1;A2=1;A1=1;A0=1;B3=0;B2=0;B1=1;B0=0;
        #5 A3=1;A2=1;A1=1;A0=1;B3=0;B2=0;B1=1;B0=1;
        #5 A3=1;A2=1;A1=1;A0=1;B3=0;B2=1;B1=0;B0=0;
        #5 A3=1;A2=1;A1=1;A0=1;B3=0;B2=1;B1=0;B0=1;
        #5 A3=1;A2=1;A1=1;A0=1;B3=0;B2=1;B1=1;B0=0;
        #5 A3=1;A2=1;A1=1;A0=1;B3=0;B2=1;B1=1;B0=1;
        #5 A3=1;A2=1;A1=1;A0=1;B3=1;B2=0;B1=0;B0=0;
        #5 A3=1;A2=1;A1=1;A0=1;B3=1;B2=0;B1=0;B0=1;
        #5 A3=1;A2=1;A1=1;A0=1;B3=1;B2=0;B1=1;B0=0;
        #5 A3=1;A2=1;A1=1;A0=1;B3=1;B2=0;B1=1;B0=1;
        #5 A3=1;A2=1;A1=1;A0=1;B3=1;B2=1;B1=0;B0=0;
        #5 A3=1;A2=1;A1=1;A0=1;B3=1;B2=1;B1=0;B0=1;
        #5 A3=1;A2=1;A1=1;A0=1;B3=1;B2=1;B1=1;B0=0;
        #5 A3=1;A2=1;A1=1;A0=1;B3=1;B2=1;B1=1;B0=1;
        #5 $finish;
    end 
endmodule