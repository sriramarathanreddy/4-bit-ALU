* SPICE3 file created from adder_subtractor.ext - technology: scmos

.include TSMC_180nm.txt
.param SUPPLY = 1.8
.global Gnd
Vdd VDD Gnd 'SUPPLY'
.option scale=0.09u

VinASA3 ASA3 Gnd DC 'SUPPLY'
VinASA2 ASA2 Gnd DC 0
VinASA1 ASA1 Gnd DC 'SUPPLY'
VinASA0 ASA0 Gnd DC 'SUPPLY'

VinASB3 ASB3 Gnd DC 'SUPPLY'
VinASB2 ASB2 Gnd DC 'SUPPLY'
VinASB1 ASB1 Gnd DC 0
VinASB0 ASB0 Gnd DC 'SUPPLY'

VinD1 D1 Gnd PULSE('SUPPLY' 0 0ns 100ps 100ps 5n 10n)

M1000 xorB2not xorB2 VDD VDD CMOSP w=20 l=2
+  ad=220 pd=62 as=11660 ps=3286
M1001 C1 FA2S1 OUT_AS2 w_1557_n253# CMOSP w=20 l=2
+  ad=440 pd=124 as=440 ps=124
M1002 FA3S1not FA3S1 VDD VDD CMOSP w=20 l=2
+  ad=220 pd=62 as=0 ps=0
M1003 ASB3not ASB3 VDD VDD CMOSP w=20 l=2
+  ad=220 pd=62 as=0 ps=0
M1004 ASA1not ASA1 VDD VDD CMOSP w=20 l=2
+  ad=440 pd=124 as=0 ps=0
M1005 ASB0not ASB0 Gnd Gnd CMOSN w=20 l=4
+  ad=220 pd=62 as=10780 ps=3038
M1006 FA0C2 a_621_274# Gnd Gnd CMOSN w=20 l=4
+  ad=220 pd=62 as=0 ps=0
M1007 a_634_222# xorB0 Gnd Gnd CMOSN w=20 l=4
+  ad=440 pd=124 as=0 ps=0
M1008 Gnd FA1C2 a_1494_186# Gnd CMOSN w=20 l=4
+  ad=0 pd=0 as=440 ps=124
M1009 C2not FA3S1not OUT_AS3 w_1036_n338# CMOSP w=20 l=2
+  ad=440 pd=124 as=440 ps=124
M1010 FA0S1 xorB0 ASA0not Gnd CMOSN w=20 l=4
+  ad=420 pd=122 as=440 ps=124
M1011 OUT_AS2 FA2S1 C1not Gnd CMOSN w=20 l=4
+  ad=420 pd=122 as=440 ps=124
M1012 C a_972_n200# VDD w_1065_n167# CMOSP w=20 l=2
+  ad=220 pd=62 as=0 ps=0
M1013 a_803_274# D1 VDD w_840_268# CMOSP w=20 l=2
+  ad=440 pd=124 as=0 ps=0
M1014 a_1325_n112# FA2S1 a_1338_n164# Gnd CMOSN w=20 l=4
+  ad=220 pd=62 as=440 ps=124
M1015 xorB0not xorB0 VDD VDD CMOSP w=20 l=2
+  ad=220 pd=62 as=0 ps=0
M1016 a_1325_274# FA1S1 a_1338_222# Gnd CMOSN w=20 l=4
+  ad=220 pd=62 as=440 ps=124
M1017 a_621_n112# ASA3 a_634_n164# Gnd CMOSN w=20 l=4
+  ad=220 pd=62 as=440 ps=124
M1018 a_803_274# FA0S1 VDD w_784_268# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1019 D1not D1 Gnd Gnd CMOSN w=20 l=4
+  ad=1540 pd=434 as=0 ps=0
M1020 OUT_AS3 FA3S1not C2 Gnd CMOSN w=20 l=4
+  ad=420 pd=122 as=440 ps=124
M1021 a_1143_274# xorB1 VDD w_1180_268# CMOSP w=20 l=2
+  ad=440 pd=124 as=0 ps=0
M1022 D1 ASB0 xorB0 w_869_481# CMOSP w=20 l=2
+  ad=1100 pd=310 as=440 ps=124
M1023 ASA3not xorB3not FA3S1 w_725_n341# CMOSP w=20 l=2
+  ad=440 pd=124 as=440 ps=124
M1024 C1 a_1494_186# Gnd Gnd CMOSN w=20 l=4
+  ad=440 pd=124 as=0 ps=0
M1025 FA3C1 a_803_n112# Gnd Gnd CMOSN w=20 l=4
+  ad=220 pd=62 as=0 ps=0
M1026 OUT_AS0 FA0S1not D1 Gnd CMOSN w=20 l=4
+  ad=420 pd=122 as=1100 ps=310
M1027 xorB3 ASB3 D1not Gnd CMOSN w=20 l=4
+  ad=420 pd=122 as=0 ps=0
M1028 a_1143_274# ASA1 VDD w_1124_268# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1029 FA0S1not FA0S1 VDD VDD CMOSP w=20 l=2
+  ad=220 pd=62 as=0 ps=0
M1030 FA1S1not FA1S1 Gnd Gnd CMOSN w=20 l=4
+  ad=220 pd=62 as=0 ps=0
M1031 xorB2 ASB2 D1not Gnd CMOSN w=20 l=4
+  ad=420 pd=122 as=0 ps=0
M1032 a_983_232# FA0C1 VDD VDD CMOSP w=20 l=2
+  ad=440 pd=124 as=0 ps=0
M1033 C0 a_972_186# VDD w_1065_219# CMOSP w=20 l=2
+  ad=440 pd=124 as=0 ps=0
M1034 a_1156_n164# xorB2 Gnd Gnd CMOSN w=20 l=4
+  ad=440 pd=124 as=0 ps=0
M1035 a_1325_n112# C1 VDD w_1362_n118# CMOSP w=20 l=2
+  ad=440 pd=124 as=0 ps=0
M1036 D1not ASB3not xorB3 w_1359_396# CMOSP w=20 l=2
+  ad=1540 pd=434 as=440 ps=124
M1037 FA3S1 xorB3not ASA3 Gnd CMOSN w=20 l=4
+  ad=420 pd=122 as=220 ps=62
M1038 a_1325_n112# FA2S1 VDD w_1306_n118# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1039 a_621_n112# xorB3 VDD w_658_n118# CMOSP w=20 l=2
+  ad=440 pd=124 as=0 ps=0
M1040 D1not D1 VDD VDD CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1041 a_983_n154# FA3C1 VDD VDD CMOSP w=20 l=2
+  ad=440 pd=124 as=0 ps=0
M1042 xorB3 ASB3not D1 Gnd CMOSN w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1043 FA2S1 xorB2 ASA2not Gnd CMOSN w=20 l=4
+  ad=420 pd=122 as=440 ps=124
M1044 xorB2 ASB2not D1 Gnd CMOSN w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1045 xorB1 ASB1not D1 Gnd CMOSN w=20 l=4
+  ad=420 pd=122 as=0 ps=0
M1046 xorB0not xorB0 Gnd Gnd CMOSN w=20 l=4
+  ad=220 pd=62 as=0 ps=0
M1047 a_621_274# ASA0 VDD w_602_268# CMOSP w=20 l=2
+  ad=440 pd=124 as=0 ps=0
M1048 ASA2not ASA2 VDD VDD CMOSP w=20 l=2
+  ad=440 pd=124 as=0 ps=0
M1049 a_972_186# FA0C2 a_983_232# w_977_226# CMOSP w=20 l=2
+  ad=220 pd=62 as=0 ps=0
M1050 C0 FA1S1 OUT_AS1 w_1557_133# CMOSP w=20 l=2
+  ad=0 pd=0 as=440 ps=124
M1051 ASB2not ASB2 VDD VDD CMOSP w=20 l=2
+  ad=220 pd=62 as=0 ps=0
M1052 D1not D1 VDD VDD CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1053 a_1338_222# C0 Gnd Gnd CMOSN w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1054 FA3C1 a_803_n112# VDD w_895_n127# CMOSP w=20 l=2
+  ad=220 pd=62 as=0 ps=0
M1055 ASB1not ASB1 VDD VDD CMOSP w=20 l=2
+  ad=220 pd=62 as=0 ps=0
M1056 Gnd FA2C1 a_1494_n200# Gnd CMOSN w=20 l=4
+  ad=0 pd=0 as=440 ps=124
M1057 FA0C1 a_803_274# VDD w_895_259# CMOSP w=20 l=2
+  ad=220 pd=62 as=0 ps=0
M1058 Gnd FA3C2 a_972_n200# Gnd CMOSN w=20 l=4
+  ad=0 pd=0 as=440 ps=124
M1059 C1not C1 VDD VDD CMOSP w=20 l=2
+  ad=440 pd=124 as=0 ps=0
M1060 ASB3not ASB3 Gnd Gnd CMOSN w=20 l=4
+  ad=220 pd=62 as=0 ps=0
M1061 FA1C2 a_1143_274# VDD w_1235_259# CMOSP w=20 l=2
+  ad=220 pd=62 as=0 ps=0
M1062 FA2S1not FA2S1 VDD VDD CMOSP w=20 l=2
+  ad=220 pd=62 as=0 ps=0
M1063 ASA1not ASA1 Gnd Gnd CMOSN w=20 l=4
+  ad=440 pd=124 as=0 ps=0
M1064 Gnd FA0C2 a_972_186# Gnd CMOSN w=20 l=4
+  ad=0 pd=0 as=440 ps=124
M1065 ASA0not ASA0 VDD VDD CMOSP w=20 l=2
+  ad=440 pd=124 as=0 ps=0
M1066 a_1143_n112# ASA2 a_1156_n164# Gnd CMOSN w=20 l=4
+  ad=220 pd=62 as=0 ps=0
M1067 FA1S1 xorB1not ASA1 Gnd CMOSN w=20 l=4
+  ad=420 pd=122 as=220 ps=62
M1068 Gnd FA0C1 a_972_186# Gnd CMOSN w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1069 ASA2not xorB2not FA2S1 w_1247_n341# CMOSP w=20 l=2
+  ad=0 pd=0 as=440 ps=124
M1070 FA2C1 a_1325_n112# Gnd Gnd CMOSN w=20 l=4
+  ad=220 pd=62 as=0 ps=0
M1071 OUT_AS0 FA0S1 D1not Gnd CMOSN w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1072 ASA0not xorB0not FA0S1 w_725_45# CMOSP w=20 l=2
+  ad=0 pd=0 as=440 ps=124
M1073 xorB1 ASB1 D1not Gnd CMOSN w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1074 D1 ASB3 xorB3 w_1358_481# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1075 a_803_274# FA0S1 a_816_222# Gnd CMOSN w=20 l=4
+  ad=220 pd=62 as=440 ps=124
M1076 D1 ASB2 xorB2 w_1202_481# CMOSP w=20 l=2
+  ad=0 pd=0 as=440 ps=124
M1077 ASA1 xorB1 FA1S1 w_1246_130# CMOSP w=20 l=2
+  ad=220 pd=62 as=440 ps=124
M1078 D1not ASB2not xorB2 w_1203_396# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1079 FA2S1 xorB2not ASA2 Gnd CMOSN w=20 l=4
+  ad=0 pd=0 as=220 ps=62
M1080 a_621_n112# ASA3 VDD w_602_n118# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1081 D1not ASB1not xorB1 w_1048_396# CMOSP w=20 l=2
+  ad=0 pd=0 as=440 ps=124
M1082 a_621_274# xorB0 VDD w_658_268# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1083 xorB3not xorB3 Gnd Gnd CMOSN w=20 l=4
+  ad=220 pd=62 as=0 ps=0
M1084 a_1143_n112# xorB2 VDD w_1180_n118# CMOSP w=20 l=2
+  ad=440 pd=124 as=0 ps=0
M1085 a_1143_n112# ASA2 VDD w_1124_n118# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1086 a_1143_274# ASA1 a_1156_222# Gnd CMOSN w=20 l=4
+  ad=220 pd=62 as=440 ps=124
M1087 OUT_AS1 FA1S1not C0 Gnd CMOSN w=20 l=4
+  ad=420 pd=122 as=440 ps=124
M1088 C1not FA2S1not OUT_AS2 w_1558_n338# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1089 ASA3not ASA3 Gnd Gnd CMOSN w=20 l=4
+  ad=440 pd=124 as=0 ps=0
M1090 a_1494_n200# FA2C2 a_1505_n154# w_1499_n160# CMOSP w=20 l=2
+  ad=220 pd=62 as=440 ps=124
M1091 FA0S1not FA0S1 Gnd Gnd CMOSN w=20 l=4
+  ad=220 pd=62 as=0 ps=0
M1092 C2 FA3S1 OUT_AS3 w_1035_n253# CMOSP w=20 l=2
+  ad=440 pd=124 as=0 ps=0
M1093 FA1C1 a_1325_274# Gnd Gnd CMOSN w=20 l=4
+  ad=220 pd=62 as=0 ps=0
M1094 FA2C1 a_1325_n112# VDD w_1417_n127# CMOSP w=20 l=2
+  ad=220 pd=62 as=0 ps=0
M1095 a_1505_232# FA1C1 VDD VDD CMOSP w=20 l=2
+  ad=440 pd=124 as=0 ps=0
M1096 D1 FA0S1 OUT_AS0 w_1035_133# CMOSP w=20 l=2
+  ad=0 pd=0 as=440 ps=124
M1097 C2not C2 Gnd Gnd CMOSN w=20 l=4
+  ad=440 pd=124 as=0 ps=0
M1098 OUT_AS2 FA2S1not C1 Gnd CMOSN w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1099 FA3C2 a_621_n112# VDD w_713_n127# CMOSP w=20 l=2
+  ad=220 pd=62 as=0 ps=0
M1100 xorB0 ASB0 D1not Gnd CMOSN w=20 l=4
+  ad=420 pd=122 as=0 ps=0
M1101 D1not FA0S1not OUT_AS0 w_1036_48# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1102 C1 a_1494_186# VDD w_1587_219# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1103 FA3S1not FA3S1 Gnd Gnd CMOSN w=20 l=4
+  ad=220 pd=62 as=0 ps=0
M1104 xorB3not xorB3 VDD VDD CMOSP w=20 l=2
+  ad=220 pd=62 as=0 ps=0
M1105 ASB2not ASB2 Gnd Gnd CMOSN w=20 l=4
+  ad=220 pd=62 as=0 ps=0
M1106 ASA3 xorB3 FA3S1 w_724_n256# CMOSP w=20 l=2
+  ad=220 pd=62 as=0 ps=0
M1107 a_816_n164# C2 Gnd Gnd CMOSN w=20 l=4
+  ad=440 pd=124 as=0 ps=0
M1108 ASB1not ASB1 Gnd Gnd CMOSN w=20 l=4
+  ad=220 pd=62 as=0 ps=0
M1109 a_816_222# D1 Gnd Gnd CMOSN w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1110 a_1494_186# FA1C2 a_1505_232# w_1499_226# CMOSP w=20 l=2
+  ad=220 pd=62 as=0 ps=0
M1111 xorB0 ASB0not D1 Gnd CMOSN w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1112 xorB1not xorB1 Gnd Gnd CMOSN w=20 l=4
+  ad=220 pd=62 as=0 ps=0
M1113 a_1156_222# xorB1 Gnd Gnd CMOSN w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1114 Gnd FA3C1 a_972_n200# Gnd CMOSN w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1115 FA3C2 a_621_n112# Gnd Gnd CMOSN w=20 l=4
+  ad=220 pd=62 as=0 ps=0
M1116 ASB0not ASB0 VDD VDD CMOSP w=20 l=2
+  ad=220 pd=62 as=0 ps=0
M1117 FA0C2 a_621_274# VDD w_713_259# CMOSP w=20 l=2
+  ad=220 pd=62 as=0 ps=0
M1118 FA2C2 a_1143_n112# Gnd Gnd CMOSN w=20 l=4
+  ad=220 pd=62 as=0 ps=0
M1119 ASA0not ASA0 Gnd Gnd CMOSN w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1120 C0 a_972_186# Gnd Gnd CMOSN w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1121 a_1325_274# C0 VDD w_1362_268# CMOSP w=20 l=2
+  ad=440 pd=124 as=0 ps=0
M1122 C2 a_1494_n200# Gnd Gnd CMOSN w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1123 D1 ASB1 xorB1 w_1047_481# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1124 xorB2not xorB2 Gnd Gnd CMOSN w=20 l=4
+  ad=220 pd=62 as=0 ps=0
M1125 xorB1not xorB1 VDD VDD CMOSP w=20 l=2
+  ad=220 pd=62 as=0 ps=0
M1126 a_1325_274# FA1S1 VDD w_1306_268# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1127 C0not C0 Gnd Gnd CMOSN w=20 l=4
+  ad=440 pd=124 as=0 ps=0
M1128 ASA2not ASA2 Gnd Gnd CMOSN w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1129 Gnd FA2C2 a_1494_n200# Gnd CMOSN w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1130 Gnd FA1C1 a_1494_186# Gnd CMOSN w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1131 a_803_n112# FA3S1 a_816_n164# Gnd CMOSN w=20 l=4
+  ad=220 pd=62 as=0 ps=0
M1132 ASA0 xorB0 FA0S1 w_724_130# CMOSP w=20 l=2
+  ad=220 pd=62 as=0 ps=0
M1133 FA1S1not FA1S1 VDD VDD CMOSP w=20 l=2
+  ad=220 pd=62 as=0 ps=0
M1134 a_1505_n154# FA2C1 VDD VDD CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1135 a_621_274# ASA0 a_634_222# Gnd CMOSN w=20 l=4
+  ad=220 pd=62 as=0 ps=0
M1136 FA2C2 a_1143_n112# VDD w_1235_n127# CMOSP w=20 l=2
+  ad=220 pd=62 as=0 ps=0
M1137 C0not C0 VDD VDD CMOSP w=20 l=2
+  ad=440 pd=124 as=0 ps=0
M1138 ASA1not xorB1not FA1S1 w_1247_45# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1139 D1not D1 Gnd Gnd CMOSN w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1140 OUT_AS3 FA3S1 C2not Gnd CMOSN w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1141 C2 a_1494_n200# VDD w_1587_n167# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1142 D1not ASB0not xorB0 w_870_396# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1143 ASA3not ASA3 VDD VDD CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1144 a_1338_n164# C1 Gnd Gnd CMOSN w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1145 FA0C1 a_803_274# Gnd Gnd CMOSN w=20 l=4
+  ad=220 pd=62 as=0 ps=0
M1146 ASA2 xorB2 FA2S1 w_1246_n256# CMOSP w=20 l=2
+  ad=220 pd=62 as=0 ps=0
M1147 a_972_n200# FA3C2 a_983_n154# w_977_n160# CMOSP w=20 l=2
+  ad=220 pd=62 as=0 ps=0
M1148 a_634_n164# xorB3 Gnd Gnd CMOSN w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1149 a_803_n112# C2 VDD w_840_n118# CMOSP w=20 l=2
+  ad=440 pd=124 as=0 ps=0
M1150 a_803_n112# FA3S1 VDD w_784_n118# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1151 C a_972_n200# Gnd Gnd CMOSN w=20 l=4
+  ad=220 pd=62 as=0 ps=0
M1152 C1not C1 Gnd Gnd CMOSN w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1153 FA1C2 a_1143_274# Gnd Gnd CMOSN w=20 l=4
+  ad=220 pd=62 as=0 ps=0
M1154 FA3S1 xorB3 ASA3not Gnd CMOSN w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1155 C0not FA1S1not OUT_AS1 w_1558_48# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1156 FA1C1 a_1325_274# VDD w_1417_259# CMOSP w=20 l=2
+  ad=220 pd=62 as=0 ps=0
M1157 OUT_AS1 FA1S1 C0not Gnd CMOSN w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1158 FA0S1 xorB0not ASA0 Gnd CMOSN w=20 l=4
+  ad=0 pd=0 as=220 ps=62
M1159 C2not C2 VDD VDD CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1160 FA2S1not FA2S1 Gnd Gnd CMOSN w=20 l=4
+  ad=220 pd=62 as=0 ps=0
M1161 FA1S1 xorB1 ASA1not Gnd CMOSN w=20 l=4
+  ad=0 pd=0 as=0 ps=0
C0 FA3S1 w_725_n341# 0.09fF
C1 w_1358_481# xorB3 0.09fF
C2 a_1494_n200# FA2C2 0.25fF
C3 FA2C2 w_1499_n160# 0.06fF
C4 w_1124_n118# VDD 0.06fF
C5 w_658_n118# VDD 0.06fF
C6 OUT_AS0 D1not 0.68fF
C7 a_803_n112# VDD 0.41fF
C8 Gnd a_634_n164# 0.21fF
C9 Gnd VDD 4.12fF
C10 VDD ASA3not 0.34fF
C11 w_1499_226# a_1494_186# 0.06fF
C12 w_1557_133# FA1S1 0.06fF
C13 w_1558_n338# FA2S1not 0.06fF
C14 VDD FA1C2 0.21fF
C15 w_724_130# ASA0 0.06fF
C16 w_1235_259# FA1C2 0.06fF
C17 w_869_481# xorB0 0.09fF
C18 w_840_268# VDD 0.06fF
C19 a_1338_n164# a_1325_n112# 0.21fF
C20 FA0S1 a_803_274# 0.29fF
C21 w_1359_396# ASB3not 0.06fF
C22 a_1143_274# a_1156_222# 0.21fF
C23 VDD a_983_232# 0.34fF
C24 w_1180_268# a_1143_274# 0.06fF
C25 w_1499_226# a_1505_232# 0.09fF
C26 w_658_268# a_621_274# 0.06fF
C27 FA3C1 Gnd 0.36fF
C28 xorB2 D1not 0.68fF
C29 ASA2 a_1143_n112# 0.29fF
C30 Gnd OUT_AS0 0.60fF
C31 w_1180_268# VDD 0.06fF
C32 FA0S1 xorB0not 0.25fF
C33 xorB0 ASA0not 0.04fF
C34 FA1S1 xorB1not 0.25fF
C35 FA2C2 w_1235_n127# 0.06fF
C36 w_724_n256# FA3S1 0.09fF
C37 a_634_222# a_621_274# 0.21fF
C38 w_1065_n167# C 0.06fF
C39 VDD ASB0 0.06fF
C40 w_1035_n253# C2 0.06fF
C41 w_1048_396# D1not 0.06fF
C42 w_977_n160# a_972_n200# 0.06fF
C43 w_1047_481# ASB1 0.06fF
C44 w_1558_48# C0not 0.06fF
C45 w_658_n118# a_621_n112# 0.06fF
C46 VDD FA0S1not 0.34fF
C47 FA1S1not Gnd 0.21fF
C48 FA1S1not OUT_AS1 0.25fF
C49 FA3S1 FA3S1not 0.04fF
C50 Gnd xorB3not 0.21fF
C51 C2 OUT_AS3 0.68fF
C52 w_1235_n127# a_1143_n112# 0.06fF
C53 Gnd FA2S1not 0.21fF
C54 FA2S1 ASA2not 0.68fF
C55 a_803_274# D1 0.16fF
C56 Gnd FA1C1 0.36fF
C57 xorB3 w_1359_396# 0.09fF
C58 w_1036_n338# OUT_AS3 0.09fF
C59 xorB0 w_658_268# 0.06fF
C60 FA0S1not OUT_AS0 0.25fF
C61 Gnd a_972_186# 0.41fF
C62 FA3S1 VDD 0.06fF
C63 ASA1not VDD 0.34fF
C64 w_1362_n118# C1 0.06fF
C65 VDD C1 0.27fF
C66 a_1494_186# a_1505_232# 0.27fF
C67 FA1S1 VDD 0.06fF
C68 w_1246_130# xorB1 0.06fF
C69 ASA3 w_724_n256# 0.06fF
C70 VDD ASA2not 0.34fF
C71 VDD FA0C2 0.21fF
C72 Gnd ASB3not 0.21fF
C73 w_713_259# VDD 0.06fF
C74 xorB0 ASB0not 0.25fF
C75 xorB0 a_621_274# 0.16fF
C76 a_1494_n200# Gnd 0.41fF
C77 ASA2 w_1124_n118# 0.06fF
C78 w_977_n160# a_983_n154# 0.09fF
C79 w_1203_396# ASB2not 0.06fF
C80 a_983_232# a_972_186# 0.27fF
C81 w_1417_259# a_1325_274# 0.06fF
C82 xorB3 D1not 0.68fF
C83 Gnd ASA0not 0.21fF
C84 w_895_259# a_803_274# 0.06fF
C85 xorB1 D1not 0.68fF
C86 VDD ASB2not 0.34fF
C87 VDD ASB1not 0.34fF
C88 VDD a_803_274# 0.41fF
C89 w_1035_n253# OUT_AS3 0.09fF
C90 a_1325_274# C0 0.16fF
C91 w_869_481# ASB0 0.06fF
C92 w_658_n118# xorB3 0.06fF
C93 w_1558_48# FA1S1not 0.06fF
C94 ASB1not ASB1 0.04fF
C95 w_895_n127# a_803_n112# 0.06fF
C96 VDD xorB0not 0.34fF
C97 w_1180_n118# a_1143_n112# 0.06fF
C98 ASA3 VDD 0.06fF
C99 a_803_n112# C2 0.16fF
C100 w_1557_n253# C1 0.06fF
C101 w_1036_48# OUT_AS0 0.09fF
C102 FA3S1 xorB3not 0.25fF
C103 Gnd C2 0.14fF
C104 xorB3 ASA3not 0.04fF
C105 FA2C1 w_1417_n127# 0.06fF
C106 FA1S1not FA1S1 0.04fF
C107 Gnd xorB2not 0.21fF
C108 xorB2 ASA2not 0.04fF
C109 Gnd FA0C1 0.36fF
C110 FA3S1not C2not 0.01fF
C111 w_1247_45# ASA1not 0.06fF
C112 w_1247_45# FA1S1 0.09fF
C113 FA0S1 ASA0 0.68fF
C114 w_602_268# ASA0 0.06fF
C115 w_840_n118# VDD 0.06fF
C116 a_1156_n164# a_1143_n112# 0.21fF
C117 Gnd a_634_222# 0.21fF
C118 w_1247_n341# ASA2not 0.06fF
C119 OUT_AS2 w_1558_n338# 0.09fF
C120 C1not VDD 0.34fF
C121 a_983_n154# a_972_n200# 0.27fF
C122 FA0C1 a_983_232# 0.05fF
C123 a_1338_222# a_1325_274# 0.21fF
C124 Gnd C 0.14fF
C125 w_1587_219# C1 0.06fF
C126 FA0S1 VDD 0.06fF
C127 xorB1 w_1180_268# 0.06fF
C128 VDD C2not 0.34fF
C129 w_1035_133# FA0S1 0.06fF
C130 FA0C2 a_972_186# 0.25fF
C131 a_1338_n164# Gnd 0.21fF
C132 xorB2 ASB2not 0.25fF
C133 Gnd ASB0not 0.21fF
C134 w_602_268# VDD 0.06fF
C135 w_1246_130# ASA1 0.06fF
C136 w_1047_481# xorB1 0.09fF
C137 ASA3 w_602_n118# 0.06fF
C138 VDD a_1505_232# 0.34fF
C139 w_1048_396# ASB1not 0.06fF
C140 w_1306_268# a_1325_274# 0.06fF
C141 w_784_268# a_803_274# 0.06fF
C142 Gnd C0 0.14fF
C143 OUT_AS1 C0 0.68fF
C144 FA2C2 Gnd 0.42fF
C145 w_977_226# a_972_186# 0.06fF
C146 w_1362_268# VDD 0.06fF
C147 xorB0 D1not 0.68fF
C148 ASA3 a_621_n112# 0.29fF
C149 w_1417_n127# VDD 0.06fF
C150 w_1359_396# D1not 0.06fF
C151 VDD ASB3 0.06fF
C152 w_1124_n118# a_1143_n112# 0.06fF
C153 ASB0not ASB0 0.04fF
C154 w_784_n118# a_803_n112# 0.06fF
C155 VDD D1 0.13fF
C156 w_1035_133# D1 0.06fF
C157 FA2C1 VDD 0.27fF
C158 OUT_AS2 Gnd 0.60fF
C159 VDD xorB1not 0.34fF
C160 ASA1not xorB1 0.04fF
C161 C1not FA2S1not 0.01fF
C162 Gnd OUT_AS3 0.60fF
C163 w_1202_481# D1 0.06fF
C164 Gnd a_1338_222# 0.21fF
C165 w_725_n341# xorB3not 0.06fF
C166 a_1325_n112# C1 0.16fF
C167 FA0S1 w_784_268# 0.06fF
C168 w_713_n127# VDD 0.06fF
C169 D1 OUT_AS0 0.68fF
C170 a_1156_n164# Gnd 0.21fF
C171 a_983_n154# VDD 0.34fF
C172 a_803_n112# a_816_n164# 0.21fF
C173 Gnd a_816_n164# 0.21fF
C174 FA2S1 VDD 0.06fF
C175 C0not VDD 0.34fF
C176 w_724_130# xorB0 0.06fF
C177 VDD FA3S1not 0.34fF
C178 FA1C1 a_1505_232# 0.05fF
C179 w_1587_219# a_1494_186# 0.06fF
C180 VDD ASA0 0.06fF
C181 w_895_259# VDD 0.06fF
C182 xorB1 ASB1not 0.25fF
C183 VDD a_1143_274# 0.41fF
C184 w_870_396# ASB0not 0.06fF
C185 w_1235_259# a_1143_274# 0.06fF
C186 xorB2 D1 0.68fF
C187 FA3C1 a_983_n154# 0.05fF
C188 w_713_259# a_621_274# 0.06fF
C189 FA3C2 Gnd 0.42fF
C190 w_1362_n118# VDD 0.06fF
C191 Gnd D1not 0.41fF
C192 w_1235_259# VDD 0.06fF
C193 FA0S1 ASA0not 0.68fF
C194 w_1035_n253# FA3S1 0.06fF
C195 w_1247_45# xorB1not 0.06fF
C196 VDD ASB1 0.06fF
C197 w_1124_268# a_1143_274# 0.06fF
C198 FA2C1 a_1505_n154# 0.05fF
C199 w_1124_268# VDD 0.06fF
C200 ASB3not ASB3 0.04fF
C201 w_784_n118# FA3S1 0.06fF
C202 w_840_n118# C2 0.06fF
C203 FA3C1 VDD 0.27fF
C204 w_1587_n167# VDD 0.06fF
C205 w_713_n127# a_621_n112# 0.06fF
C206 w_725_45# xorB0not 0.06fF
C207 w_1035_133# OUT_AS0 0.09fF
C208 w_1557_n253# FA2S1 0.06fF
C209 OUT_AS2 C1 0.68fF
C210 OUT_AS1 Gnd 0.60fF
C211 FA1S1not C0not 0.01fF
C212 Gnd ASA3not 0.21fF
C213 w_869_481# D1 0.06fF
C214 FA2S1 FA2S1not 0.04fF
C215 xorB2 w_1203_396# 0.09fF
C216 Gnd FA1C2 0.42fF
C217 w_1036_n338# C2not 0.06fF
C218 FA1S1 ASA1 0.68fF
C219 w_870_396# xorB0 0.09fF
C220 w_1306_n118# FA2S1 0.06fF
C221 w_602_n118# VDD 0.06fF
C222 FA2S1 w_1247_n341# 0.09fF
C223 FA0S1not D1not 0.01fF
C224 Gnd a_1156_222# 0.21fF
C225 FA1S1 a_1325_274# 0.29fF
C226 xorB2 VDD 0.06fF
C227 FA1S1not VDD 0.34fF
C228 VDD xorB3not 0.34fF
C229 a_621_n112# VDD 0.41fF
C230 a_621_n112# a_634_n164# 0.21fF
C231 FA1S1 w_1306_268# 0.06fF
C232 w_1246_130# FA1S1 0.09fF
C233 w_725_45# FA0S1 0.09fF
C234 VDD FA2S1not 0.34fF
C235 VDD FA1C1 0.27fF
C236 w_1202_481# xorB2 0.09fF
C237 w_784_268# VDD 0.06fF
C238 w_1306_n118# VDD 0.06fF
C239 w_1417_n127# a_1325_n112# 0.06fF
C240 a_1505_n154# VDD 0.34fF
C241 xorB3 D1 0.68fF
C242 w_602_268# a_621_274# 0.06fF
C243 w_1358_481# ASB3 0.06fF
C244 Gnd FA0S1not 0.21fF
C245 w_1587_219# VDD 0.06fF
C246 xorB1 D1 0.68fF
C247 ASA2 FA2S1 0.68fF
C248 w_1065_219# VDD 0.06fF
C249 w_724_n256# xorB3 0.06fF
C250 w_1358_481# D1 0.06fF
C251 w_1065_n167# a_972_n200# 0.06fF
C252 VDD ASB3not 0.34fF
C253 w_870_396# D1not 0.06fF
C254 w_1246_n256# FA2S1 0.09fF
C255 ASB2not ASB2 0.04fF
C256 w_1558_48# OUT_AS1 0.09fF
C257 OUT_AS2 C1not 0.68fF
C258 w_602_n118# a_621_n112# 0.06fF
C259 VDD ASA0not 0.34fF
C260 w_1362_268# C0 0.06fF
C261 w_1557_133# C0 0.06fF
C262 ASA2 VDD 0.06fF
C263 FA3S1 a_803_n112# 0.29fF
C264 FA3S1 Gnd 0.31fF
C265 ASA1not Gnd 0.21fF
C266 w_1036_48# D1not 0.06fF
C267 FA3S1 ASA3not 0.68fF
C268 Gnd C1 0.14fF
C269 FA1S1 Gnd 0.31fF
C270 FA2S1 xorB2not 0.25fF
C271 Gnd ASA2not 0.21fF
C272 Gnd FA0C2 0.42fF
C273 OUT_AS3 C2not 0.68fF
C274 FA2S1 a_1325_n112# 0.29fF
C275 a_1494_n200# w_1587_n167# 0.06fF
C276 w_1036_n338# FA3S1not 0.06fF
C277 FA3C2 w_977_n160# 0.06fF
C278 w_895_259# FA0C1 0.06fF
C279 w_895_n127# VDD 0.06fF
C280 Gnd a_816_222# 0.21fF
C281 xorB1 a_1143_274# 0.16fF
C282 C1not w_1558_n338# 0.06fF
C283 xorB3 VDD 0.06fF
C284 VDD C2 0.27fF
C285 xorB1 VDD 0.06fF
C286 VDD xorB2not 0.34fF
C287 w_1235_n127# VDD 0.06fF
C288 w_1362_n118# a_1325_n112# 0.06fF
C289 VDD FA0C1 0.27fF
C290 w_1499_226# FA1C2 0.06fF
C291 a_1325_n112# VDD 0.41fF
C292 Gnd ASB2not 0.21fF
C293 w_658_268# VDD 0.06fF
C294 Gnd ASB1not 0.21fF
C295 FA3C1 w_895_n127# 0.06fF
C296 ASA0 a_621_274# 0.29fF
C297 w_1362_268# a_1325_274# 0.06fF
C298 w_977_226# a_983_232# 0.09fF
C299 w_840_268# a_803_274# 0.06fF
C300 Gnd xorB0not 0.21fF
C301 xorB0 D1 0.68fF
C302 w_1587_n167# C2 0.06fF
C303 w_1065_219# a_972_186# 0.06fF
C304 C VDD 0.21fF
C305 w_1417_259# VDD 0.06fF
C306 a_1494_n200# a_1505_n154# 0.27fF
C307 w_1065_n167# VDD 0.06fF
C308 w_1499_n160# a_1505_n154# 0.09fF
C309 VDD ASB0not 0.34fF
C310 VDD a_621_274# 0.41fF
C311 w_1246_n256# xorB2 0.06fF
C312 w_840_n118# a_803_n112# 0.06fF
C313 VDD C0 0.27fF
C314 FA2C2 VDD 0.21fF
C315 FA3C2 a_972_n200# 0.25fF
C316 C1not Gnd 0.21fF
C317 w_1036_48# FA0S1not 0.06fF
C318 a_1494_n200# w_1499_n160# 0.06fF
C319 FA0S1 Gnd 0.31fF
C320 a_621_n112# xorB3 0.16fF
C321 ASA1not FA1S1 0.68fF
C322 Gnd C2not 0.21fF
C323 Gnd a_1494_186# 0.41fF
C324 FA3S1not OUT_AS3 0.25fF
C325 w_725_n341# ASA3not 0.06fF
C326 a_1494_186# FA1C2 0.25fF
C327 w_1048_396# xorB1 0.09fF
C328 w_713_259# FA0C2 0.06fF
C329 w_784_n118# VDD 0.06fF
C330 w_1247_n341# xorB2not 0.06fF
C331 w_1306_n118# a_1325_n112# 0.06fF
C332 w_1180_n118# VDD 0.06fF
C333 a_1143_n112# VDD 0.41fF
C334 Gnd a_972_n200# 0.41fF
C335 xorB0 VDD 0.06fF
C336 w_1557_133# OUT_AS1 0.09fF
C337 w_724_130# FA0S1 0.09fF
C338 ASA1 a_1143_274# 0.29fF
C339 xorB3 ASB3not 0.25fF
C340 VDD ASA1 0.06fF
C341 w_1417_259# FA1C1 0.06fF
C342 w_977_226# FA0C2 0.06fF
C343 ASA2 w_1246_n256# 0.06fF
C344 FA3C2 w_713_n127# 0.06fF
C345 VDD a_1325_274# 0.41fF
C346 ASA3 FA3S1 0.68fF
C347 FA2C1 Gnd 0.36fF
C348 w_1124_268# ASA1 0.06fF
C349 Gnd xorB1not 0.21fF
C350 w_1306_268# VDD 0.06fF
C351 FA0S1 FA0S1not 0.04fF
C352 w_840_268# D1 0.06fF
C353 w_1203_396# D1not 0.06fF
C354 a_816_222# a_803_274# 0.21fF
C355 VDD ASB2 0.06fF
C356 w_1202_481# ASB2 0.06fF
C357 w_1557_n253# OUT_AS2 0.09fF
C358 FA3C2 VDD 0.21fF
C359 w_1180_n118# xorB2 0.06fF
C360 VDD D1not 0.67fF
C361 w_1065_219# C0 0.06fF
C362 w_725_45# ASA0not 0.06fF
C363 xorB2 a_1143_n112# 0.16fF
C364 Gnd FA2S1 0.31fF
C365 C0not Gnd 0.21fF
C366 OUT_AS1 C0not 0.68fF
C367 Gnd FA3S1not 0.21fF
C368 OUT_AS2 FA2S1not 0.25fF
C369 w_1047_481# D1 0.06fF
C370 FA2S1 Gnd 1.27fF
C371 Gnd Gnd 1.75fF
C372 xorB2 Gnd 1.30fF
C373 FA3S1 Gnd 1.75fF
C374 xorB3 Gnd 1.58fF
C375 C1not Gnd 0.22fF
C376 OUT_AS2 Gnd 0.03fF
C377 FA2S1not Gnd 0.54fF
C378 ASA2not Gnd 0.24fF
C379 xorB2not Gnd 0.62fF
C380 C2not Gnd 0.02fF
C381 OUT_AS3 Gnd 0.78fF
C382 FA3S1not Gnd 0.43fF
C383 ASA3not Gnd 0.13fF
C384 xorB3not Gnd 0.53fF
C385 C1 Gnd 0.53fF
C386 C2 Gnd 0.73fF
C387 ASA2 Gnd 0.55fF
C388 ASA3 Gnd 0.85fF
C389 FA2C2 Gnd 0.45fF
C390 FA2C1 Gnd 0.14fF
C391 FA3C2 Gnd 0.46fF
C392 FA3C1 Gnd 0.46fF
C393 a_1494_n200# Gnd 0.77fF
C394 a_1338_n164# Gnd 0.18fF
C395 a_1156_n164# Gnd 0.18fF
C396 C Gnd 0.13fF
C397 a_972_n200# Gnd 0.77fF
C398 a_816_n164# Gnd 0.18fF
C399 a_634_n164# Gnd 0.18fF
C400 a_1505_n154# Gnd 0.13fF
C401 a_1325_n112# Gnd 0.80fF
C402 a_1143_n112# Gnd 0.80fF
C403 a_983_n154# Gnd 0.13fF
C404 a_803_n112# Gnd 0.80fF
C405 a_621_n112# Gnd 0.80fF
C406 FA1S1 Gnd 1.15fF
C407 xorB1 Gnd 0.99fF
C408 FA0S1 Gnd 1.47fF
C409 xorB0 Gnd 1.66fF
C410 C0not Gnd 0.21fF
C411 OUT_AS1 Gnd 0.03fF
C412 FA1S1not Gnd 0.54fF
C413 ASA1not Gnd 0.20fF
C414 xorB1not Gnd 0.64fF
C415 D1not Gnd 0.59fF
C416 OUT_AS0 Gnd 0.77fF
C417 FA0S1not Gnd 0.43fF
C418 ASA0not Gnd 0.11fF
C419 xorB0not Gnd 0.54fF
C420 C0 Gnd 0.72fF
C421 D1 Gnd 1.18fF
C422 ASA1 Gnd 0.54fF
C423 ASA0 Gnd 0.78fF
C424 FA1C2 Gnd 0.42fF
C425 FA1C1 Gnd 0.14fF
C426 FA0C2 Gnd 0.43fF
C427 FA0C1 Gnd 0.46fF
C428 a_1494_186# Gnd 0.77fF
C429 a_1338_222# Gnd 0.22fF
C430 a_1156_222# Gnd 0.11fF
C431 a_972_186# Gnd 0.77fF
C432 a_816_222# Gnd 0.22fF
C433 a_634_222# Gnd 0.22fF
C434 a_1505_232# Gnd 0.13fF
C435 a_1325_274# Gnd 0.39fF
C436 a_1143_274# Gnd 0.33fF
C437 a_983_232# Gnd 0.13fF
C438 a_803_274# Gnd 0.44fF
C439 a_621_274# Gnd 0.41fF
C440 ASB3 Gnd 0.38fF
C441 ASB2 Gnd 0.85fF
C442 ASB1 Gnd 0.64fF
C443 ASB0 Gnd 0.53fF
C444 ASB3not Gnd 0.54fF
C445 ASB2not Gnd 0.66fF
C446 ASB1not Gnd 0.66fF
C447 ASB0not Gnd 0.33fF
C448 w_1558_n338# Gnd 0.93fF
C449 VDD Gnd 17.55fF
C450 w_1247_n341# Gnd 1.16fF
C451 w_1036_n338# Gnd 1.16fF
C452 w_725_n341# Gnd 1.16fF
C453 w_1557_n253# Gnd 0.96fF
C454 w_1246_n256# Gnd 1.16fF
C455 w_1035_n253# Gnd 1.16fF
C456 w_724_n256# Gnd 1.16fF
C457 w_1587_n167# Gnd 1.16fF
C458 w_1499_n160# Gnd 0.13fF
C459 w_1065_n167# Gnd 1.16fF
C460 w_977_n160# Gnd 0.13fF
C461 w_1417_n127# Gnd 1.16fF
C462 w_1362_n118# Gnd 1.16fF
C463 w_1306_n118# Gnd 1.16fF
C464 w_1235_n127# Gnd 1.16fF
C465 w_1180_n118# Gnd 1.16fF
C466 w_1124_n118# Gnd 1.16fF
C467 w_895_n127# Gnd 1.16fF
C468 w_840_n118# Gnd 1.16fF
C469 w_784_n118# Gnd 1.16fF
C470 w_713_n127# Gnd 1.16fF
C471 w_658_n118# Gnd 1.16fF
C472 w_602_n118# Gnd 1.16fF
C473 w_1558_48# Gnd 0.93fF
C474 w_1247_45# Gnd 1.16fF
C475 w_1036_48# Gnd 1.16fF
C476 w_725_45# Gnd 1.16fF
C477 w_1557_133# Gnd 0.96fF
C478 w_1246_130# Gnd 1.16fF
C479 w_1035_133# Gnd 1.16fF
C480 w_724_130# Gnd 1.16fF
C481 w_1587_219# Gnd 1.16fF
C482 w_1499_226# Gnd 0.13fF
C483 w_1065_219# Gnd 1.16fF
C484 w_977_226# Gnd 0.13fF
C485 w_1417_259# Gnd 1.16fF
C486 w_1362_268# Gnd 0.80fF
C487 w_1306_268# Gnd 1.16fF
C488 w_1235_259# Gnd 1.16fF
C489 w_1180_268# Gnd 0.00fF
C490 w_1124_268# Gnd 1.16fF
C491 w_840_268# Gnd 1.16fF
C492 w_713_259# Gnd 1.16fF
C493 w_658_268# Gnd 0.93fF
C494 w_602_268# Gnd 1.16fF
C495 w_1359_396# Gnd 0.17fF
C496 w_1203_396# Gnd 0.61fF
C497 w_1048_396# Gnd 0.61fF
C498 w_870_396# Gnd 1.16fF
C499 w_1358_481# Gnd 0.93fF
C500 w_1202_481# Gnd 1.16fF
C501 w_1047_481# Gnd 1.16fF
C502 w_869_481# Gnd 0.58fF

.tran 1n 10n
.control
run
set color0 = white
set color1 = black
plot v(OUT_AS0) v(OUT_AS1)+2 v(OUT_AS2)+4 v(OUT_AS3)+6 v(C)+8 v(D1)+10
.endc
.end