magic
tech scmos
timestamp 1701785186
<< nwell >>
rect 415 58 437 86
rect 533 83 555 111
rect 485 54 507 82
rect 556 4 578 32
<< ntransistor >>
rect 562 95 572 99
rect 421 39 431 43
rect 491 35 501 39
rect 539 16 549 20
<< ptransistor >>
rect 539 96 549 98
rect 421 71 431 73
rect 491 67 501 69
rect 562 17 572 19
<< ndiffusion >>
rect 562 99 572 100
rect 562 94 572 95
rect 421 43 431 44
rect 491 39 501 40
rect 421 38 431 39
rect 491 34 501 35
rect 539 20 549 21
rect 539 15 549 16
<< pdiffusion >>
rect 539 98 549 100
rect 539 94 549 96
rect 421 73 431 75
rect 421 69 431 71
rect 491 69 501 71
rect 491 65 501 67
rect 562 19 572 21
rect 562 15 572 17
<< ndcontact >>
rect 562 100 572 105
rect 562 89 572 94
rect 421 44 431 49
rect 491 40 501 45
rect 421 33 431 38
rect 491 29 501 34
rect 539 21 549 26
rect 539 10 549 15
<< pdcontact >>
rect 539 100 549 105
rect 539 89 549 94
rect 421 75 431 80
rect 491 71 501 76
rect 421 64 431 69
rect 491 60 501 65
rect 562 21 572 26
rect 562 10 572 15
<< psubstratepcontact >>
rect 424 25 428 29
rect 494 21 498 25
<< nsubstratencontact >>
rect 542 111 546 116
rect 424 86 428 90
rect 494 82 498 86
rect 565 32 569 36
<< polysilicon >>
rect 450 98 527 100
rect 522 96 539 98
rect 549 96 552 98
rect 559 95 562 99
rect 572 98 575 99
rect 572 96 584 98
rect 572 95 575 96
rect 437 86 475 90
rect 471 82 485 86
rect 413 71 421 73
rect 431 71 434 73
rect 483 67 491 69
rect 501 67 504 69
rect 511 52 515 89
rect 582 57 584 96
rect 582 55 592 57
rect 418 42 421 43
rect 413 40 421 42
rect 418 39 421 40
rect 431 39 434 43
rect 488 38 491 39
rect 483 36 491 38
rect 488 35 491 36
rect 501 35 504 39
rect 439 25 483 29
rect 479 21 487 25
rect 536 19 539 20
rect 450 17 475 19
rect 472 14 475 17
rect 495 17 539 19
rect 495 14 498 17
rect 536 16 539 17
rect 549 16 552 20
rect 582 19 584 55
rect 559 17 562 19
rect 572 17 584 19
rect 472 12 498 14
rect 590 3 592 55
rect 457 1 592 3
<< polycontact >>
rect 446 97 450 101
rect 433 86 437 90
rect 511 89 515 94
rect 485 82 489 86
rect 503 82 507 86
rect 409 70 413 74
rect 479 66 483 70
rect 511 48 515 52
rect 409 39 413 43
rect 479 35 483 39
rect 435 25 439 29
rect 487 21 491 25
rect 446 16 450 20
rect 453 0 457 4
<< metal1 >>
rect 538 111 542 116
rect 546 111 555 116
rect 394 97 446 101
rect 549 100 562 105
rect 572 100 610 105
rect 394 56 398 97
rect 415 86 424 90
rect 428 86 433 90
rect 515 89 539 94
rect 549 89 562 94
rect 424 80 428 86
rect 489 82 494 86
rect 498 82 503 86
rect 507 82 522 86
rect 494 76 498 82
rect 409 56 413 70
rect 389 52 413 56
rect 394 20 398 52
rect 409 43 413 52
rect 424 56 428 64
rect 479 56 483 66
rect 424 52 457 56
rect 466 52 483 56
rect 424 49 428 52
rect 424 29 428 33
rect 421 25 424 29
rect 428 25 435 29
rect 394 16 446 20
rect 453 4 457 52
rect 472 10 476 52
rect 479 39 483 52
rect 494 52 498 60
rect 494 48 511 52
rect 494 45 498 48
rect 523 36 527 81
rect 606 58 610 100
rect 606 54 617 58
rect 523 32 565 36
rect 569 32 578 36
rect 494 25 498 29
rect 491 21 494 25
rect 498 21 501 25
rect 515 21 539 26
rect 549 21 562 26
rect 515 10 519 21
rect 606 15 610 54
rect 549 10 562 15
rect 572 10 610 15
rect 472 5 519 10
<< m2contact >>
rect 533 111 538 116
rect 522 81 527 86
<< metal2 >>
rect 522 111 533 116
rect 522 86 527 111
<< labels >>
rlabel metal1 421 25 431 29 1 Gnd
rlabel metal1 610 54 617 58 7 Out
rlabel metal1 389 52 394 56 3 A
rlabel metal1 466 52 471 56 1 B
rlabel metal1 533 111 555 116 5 VDD
<< end >>
