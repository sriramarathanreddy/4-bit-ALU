magic
tech scmos
timestamp 1701500891
<< nwell >>
rect 213 137 249 169
rect 269 137 305 169
rect 325 137 361 169
rect 381 137 417 169
<< ntransistor >>
rect 256 91 260 111
rect 256 51 260 71
rect 256 11 260 31
rect 256 -28 260 -8
<< ptransistor >>
rect 230 143 232 163
rect 286 143 288 163
rect 342 143 344 163
rect 398 143 400 163
<< ndiffusion >>
rect 255 91 256 111
rect 260 91 261 111
rect 255 51 256 71
rect 260 51 261 71
rect 255 11 256 31
rect 260 11 261 31
rect 255 -28 256 -8
rect 260 -28 261 -8
<< pdiffusion >>
rect 229 143 230 163
rect 232 143 233 163
rect 285 143 286 163
rect 288 143 289 163
rect 341 143 342 163
rect 344 143 345 163
rect 397 143 398 163
rect 400 143 401 163
<< ndcontact >>
rect 245 91 255 111
rect 261 91 271 111
rect 245 51 255 71
rect 261 51 271 71
rect 245 11 255 31
rect 261 11 271 31
rect 245 -28 255 -8
rect 261 -28 271 -8
<< pdcontact >>
rect 219 143 229 163
rect 233 143 243 163
rect 275 143 285 163
rect 289 143 299 163
rect 331 143 341 163
rect 345 143 355 163
rect 387 143 397 163
rect 401 143 411 163
<< psubstratepcontact >>
rect 213 -37 217 -33
rect 413 -37 417 -33
<< nsubstratencontact >>
rect 213 169 217 173
rect 413 169 417 173
<< polysilicon >>
rect 230 163 232 166
rect 286 163 288 166
rect 342 163 344 166
rect 398 163 400 166
rect 230 134 232 143
rect 286 134 288 143
rect 342 134 344 143
rect 398 134 400 143
rect 217 130 232 134
rect 273 130 288 134
rect 329 130 344 134
rect 385 130 400 134
rect 245 114 260 118
rect 256 111 260 114
rect 256 88 260 91
rect 284 78 288 130
rect 245 74 288 78
rect 256 71 260 74
rect 256 48 260 51
rect 340 38 344 130
rect 245 34 344 38
rect 256 31 260 34
rect 256 8 260 11
rect 396 -1 400 130
rect 245 -5 400 -1
rect 256 -8 260 -5
rect 256 -31 260 -28
<< polycontact >>
rect 213 130 217 134
rect 241 114 245 118
rect 241 74 245 78
rect 241 34 245 38
rect 241 -5 245 -1
<< metal1 >>
rect 217 169 413 173
rect 219 163 229 169
rect 275 163 285 169
rect 331 163 341 169
rect 387 163 397 169
rect 198 130 213 134
rect 198 118 202 130
rect 233 125 243 143
rect 289 125 299 143
rect 345 125 355 143
rect 401 125 411 143
rect 213 121 417 125
rect 198 114 241 118
rect 261 111 271 121
rect 245 85 255 91
rect 245 81 271 85
rect 226 74 241 78
rect 261 71 271 81
rect 245 45 255 51
rect 245 41 271 45
rect 226 34 241 38
rect 261 31 271 41
rect 245 6 255 11
rect 245 2 271 6
rect 226 -5 241 -1
rect 261 -8 271 2
rect 245 -33 255 -28
rect 217 -37 413 -33
<< labels >>
rlabel metal1 198 130 217 134 1 A
rlabel metal1 226 74 245 78 1 B
rlabel metal1 213 169 361 173 5 VDD
rlabel metal1 226 34 245 38 1 C
rlabel metal1 213 121 417 125 1 OUT
rlabel metal1 226 -5 245 -1 1 D
rlabel metal1 213 -37 417 -33 1 Gnd
<< end >>
